library IEEE;
use IEEE.std_logic_1164.ALL;

entity spi_master_tb is
end spi_master_tb;

