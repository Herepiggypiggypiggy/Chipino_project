configuration texture_ctrl_behaviour_cfg of texture_ctrl is
   for behaviour
   end for;
end texture_ctrl_behaviour_cfg;
