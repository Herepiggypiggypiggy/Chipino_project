library IEEE;
use IEEE.std_logic_1164.all;

entity color_ctrl_tb is
end color_ctrl_tb;

