configuration not_arduino_behaviour_cfg of not_arduino is
   for behaviour
   end for;
end not_arduino_behaviour_cfg;
