library IEEE;
use IEEE.std_logic_1164.ALL;

entity player_fsm_tb is
end player_fsm_tb;
