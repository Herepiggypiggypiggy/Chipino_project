library IEEE;
use IEEE.std_logic_1164.ALL;

entity spi_v3_tb is
end spi_v3_tb;
