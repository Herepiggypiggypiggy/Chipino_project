library IEEE;
use IEEE.std_logic_1164.ALL;

entity vga_test_tb is
end vga_test_tb;
