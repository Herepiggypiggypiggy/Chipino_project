configuration tile_ctrl_behavioural_cfg of tile_ctrl is
   for behavioural
   end for;
end tile_ctrl_behavioural_cfg;
