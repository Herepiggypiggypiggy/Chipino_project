
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of module_test is

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD1P5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL02BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL015BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD10BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFQD0BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OR3XD1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component AO31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component FA1D0BWP7T
    port(A, B, CI : in std_logic; CO, S : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component OR4XD1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component MAOI222D1BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKMUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component DFCNQD1BWP7T
    port(CDN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component EDFCND1BWP7T
    port(CDN, CP, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component AOI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component DFCND1BWP7T
    port(CDN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFXD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q, QN : out std_logic);
  end component;

  component AOI221D1BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component OA222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component OAI33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D1BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D1BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component NR3D1BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D2BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1P5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OA31D2BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component AN3D2BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component EDFKCND1BWP7T
    port(CN, CP, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component ND2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D2BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  signal FE_PHN510_map_data_9, FE_PHN509_map_data_56, FE_PHN508_stable_map_com_n_86, FE_PHN507_map_data_24, FE_PHN506_map_data_30 : std_logic;
  signal FE_PHN505_map_data_42, FE_PHN504_map_data_26, FE_PHN503_map_data_40, FE_PHN502_fsm_com_n_489, FE_PHN501_map_data_26 : std_logic;
  signal FE_PHN500_map_data_16, FE_PHN499_map_data_32, FE_PHN498_level_d_1, FE_PHN497_map_data_22, FE_PHN496_map_data_15 : std_logic;
  signal FE_PHN495_map_data_45, FE_PHN494_spi_com_n_74, FE_PHN493_map_data_25, FE_PHN492_stable_map_com_n_79, FE_PHN491_map_data_29 : std_logic;
  signal FE_PHN490_map_data_31, FE_PHN489_level_d_1, FE_PHN488_stable_map_com_n_79, FE_PHN487_fsm_com_n_489, FE_PHN486_map_data_28 : std_logic;
  signal FE_PHN485_map_data_55, FE_PHN484_map_data_47, FE_PHN483_map_data_59, FE_PHN482_map_data_30, FE_PHN481_map_data_16 : std_logic;
  signal FE_PHN480_map_data_56, FE_PHN479_spi_com_n_74, FE_PHN478_map_data_50, FE_PHN477_level_d_4, FE_PHN476_map_data_21 : std_logic;
  signal FE_PHN475_map_data_15, FE_PHN474_map_data_32, FE_PHN473_map_data_39, FE_PHN472_map_data_60, FE_PHN471_stable_map_com_n_84 : std_logic;
  signal FE_PHN470_map_data_41, FE_PHN469_map_data_45, FE_PHN468_map_data_43, FE_PHN467_map_data_22, FE_PHN466_map_data_40 : std_logic;
  signal FE_PHN465_map_data_4, FE_PHN464_map_data_24, FE_PHN463_map_data_42, FE_PHN462_spi_com_MISO_shift_42, FE_PHN461_map_data_8 : std_logic;
  signal FE_PHN460_stable_map_com_n_102, FE_PHN459_fsm_com_n_489, FE_PHN458_energy_d_7, FE_PHN457_map_data_64, FE_PHN456_fsm_com_energy_8 : std_logic;
  signal FE_PHN455_spi_com_MISO_shift_42, FE_PHN454_level_d_1, FE_PHN453_spi_com_MISO_shift_34, FE_PHN452_map_data_50, FE_PHN451_map_data_59 : std_logic;
  signal FE_PHN450_map_data_16, FE_PHN449_map_data_28, FE_PHN448_map_data_60, FE_PHN447_map_data_30, FE_PHN446_map_data_32 : std_logic;
  signal FE_PHN445_map_data_40, FE_PHN444_map_data_47, FE_PHN443_map_data_43, FE_PHN442_map_data_22, FE_PHN441_spi_com_MISO_shift_14 : std_logic;
  signal FE_PHN440_map_data_31, FE_PHN439_map_data_11, FE_PHN438_map_data_3, FE_PHN437_map_data_29, FE_PHN436_map_data_45 : std_logic;
  signal FE_PHN435_map_data_25, FE_PHN434_map_data_39, FE_PHN433_stable_map_com_n_79, FE_PHN432_map_data_24, FE_PHN431_map_data_15 : std_logic;
  signal FE_PHN430_stable_map_com_n_102, FE_PHN429_map_data_56, FE_PHN428_map_data_55, FE_PHN427_stable_map_com_n_58, FE_PHN426_map_data_42 : std_logic;
  signal FE_PHN425_map_data_9, FE_PHN424_map_data_21, FE_PHN423_map_data_26, FE_PHN422_map_data_41, FE_PHN421_spi_com_MISO_shift_18 : std_logic;
  signal FE_PHN420_spi_com_n_74, FE_PHN419_spi_com_bit_count_0, FE_PHN418_spi_com_MISO_shift_46, FE_PHN417_map_data_8, FE_PHN416_map_data_58 : std_logic;
  signal FE_PHN415_map_data_2, FE_PHN414_map_data_4, FE_PHN413_level_d_4, FE_PHN412_stable_map_com_n_84, FE_PHN411_map_data_6 : std_logic;
  signal FE_PHN410_energy_d_11, FE_PHN409_spi_com_MISO_shift_11, FE_PHN408_vga_com_texture_module_n_193, FE_PHN407_fsm_com_n_106, FE_PHN406_spi_com_n_178 : std_logic;
  signal FE_PHN405_spi_com_n_83, FE_PHN404_vga_com_texture_module_n_252, FE_PHN403_energy_d_1, FE_PHN402_energy_d_11, FE_PHN401_vga_com_vcount_2 : std_logic;
  signal FE_PHN400_energy_d_7, FE_PHN399_fsm_com_energy_8, FE_PHN398_spi_com_MISO_shift_18, FE_PHN397_fsm_com_energy_0, FE_PHN396_fsm_com_reached_high_0 : std_logic;
  signal FE_PHN395_fsm_com_energy_3, FE_PHN394_map_data_64, FE_PHN393_stable_map_com_n_84, FE_PHN392_map_data_6, FE_PHN391_vga_com_texture_module_vvis_0 : std_logic;
  signal FE_PHN390_map_data_8, FE_PHN389_map_data_2, FE_PHN388_map_data_58, FE_PHN387_map_data_62, FE_PHN386_vga_com_texture_module_n_129 : std_logic;
  signal FE_PHN385_map_data_volatile_71, FE_PHN384_map_data_4, FE_PHN383_energy_d_10, FE_PHN382_level_d_4, FE_PHN381_map_data_volatile_46 : std_logic;
  signal FE_PHN380_spi_com_MISO_shift_40, FE_PHN379_spi_com_MOSI_shift_14, FE_PHN378_map_data_volatile_37, FE_PHN377_map_data_volatile_36, FE_PHN376_spi_com_MISO_shift_12 : std_logic;
  signal FE_PHN375_spi_com_MOSI_shift_12, FE_PHN374_spi_com_bit_count_0, FE_PHN373_n_87, FE_PHN372_n_95, FE_PHN371_spi_com_SCLK_count_1 : std_logic;
  signal FE_PHN370_vga_com_texture_module_hvis_3, FE_PHN369_spi_com_MISO_shift_34, FE_PHN368_spi_com_MISO_shift_46, FE_PHN367_spi_com_MISO_shift_14, FE_PHN366_spi_com_MISO_shift_42 : std_logic;
  signal FE_PHN365_fsm_com_n_20, FE_PHN364_map_data_volatile_10, FE_PHN363_fsm_com_n_103, FE_PHN362_vga_com_texture_module_n_176, FE_PHN361_vga_com_texture_module_n_190 : std_logic;
  signal FE_PHN360_fsm_com_n_497, FE_PHN359_fsm_com_n_225, FE_PHN358_vga_com_texture_module_n_238, FE_PHN357_fsm_com_n_298, FE_PHN356_fsm_com_n_197 : std_logic;
  signal FE_PHN355_fsm_com_n_482, FE_PHN354_vga_com_texture_module_n_239, FE_PHN353_vga_com_texture_module_n_174, FE_PHN352_vga_com_texture_module_n_52, FE_PHN351_spi_com_n_254 : std_logic;
  signal FE_PHN350_stable_map_com_n_106, FE_PHN349_stable_map_com_n_130, FE_PHN348_stable_map_com_n_134, FE_PHN347_stable_map_com_n_59, FE_PHN346_stable_map_com_n_107 : std_logic;
  signal FE_PHN345_stable_map_com_n_82, FE_PHN344_vga_com_texture_module_n_240, FE_PHN343_vga_com_texture_module_n_232, FE_PHN342_vga_com_texture_module_n_254, FE_PHN341_vga_com_texture_module_n_216 : std_logic;
  signal FE_PHN340_fsm_com_n_487, FE_PHN339_vga_com_texture_module_n_249, FE_PHN338_stable_map_com_n_49, FE_PHN337_fsm_com_n_473, FE_PHN336_fsm_com_n_378 : std_logic;
  signal FE_PHN335_vga_com_texture_module_n_251, FE_PHN334_spi_com_n_45, FE_PHN333_n_144, FE_PHN332_stable_map_com_n_55, FE_PHN331_vga_com_texture_module_n_162 : std_logic;
  signal FE_PHN330_fsm_com_n_465, FE_PHN329_fsm_com_n_363, FE_PHN328_stable_map_com_n_136, FE_PHN327_vga_com_texture_module_n_253, FE_PHN326_vga_com_texture_module_n_48 : std_logic;
  signal FE_PHN325_vga_com_texture_module_n_229, FE_PHN324_spi_com_n_246, FE_PHN323_stable_map_com_n_133, FE_PHN322_spi_com_n_257, FE_PHN321_fsm_com_n_340 : std_logic;
  signal FE_PHN320_fsm_com_n_359, FE_PHN319_spi_com_n_258, FE_PHN318_vga_com_texture_module_n_248, FE_PHN317_fsm_com_n_202, FE_PHN316_fsm_com_n_491 : std_logic;
  signal FE_PHN315_spi_com_n_224, FE_PHN314_fsm_com_n_474, FE_PHN313_fsm_com_n_472, FE_PHN312_vga_com_texture_module_n_242, FE_PHN311_vga_com_texture_module_n_201 : std_logic;
  signal FE_PHN310_stable_map_com_n_126, FE_PHN309_vga_com_texture_module_n_187, FE_PHN308_fsm_com_n_380, FE_PHN307_stable_map_com_n_60, FE_PHN306_spi_com_n_243 : std_logic;
  signal FE_PHN305_stable_map_com_n_137, FE_PHN304_fsm_com_n_477, FE_PHN303_spi_com_n_55, FE_PHN302_spi_com_n_226, FE_PHN301_spi_com_n_242 : std_logic;
  signal FE_PHN300_vga_com_texture_module_n_223, FE_PHN299_fsm_com_n_357, FE_PHN298_vga_com_texture_module_n_202, FE_PHN297_stable_map_com_n_109, FE_PHN296_fsm_com_n_464 : std_logic;
  signal FE_PHN295_spi_com_n_229, FE_PHN294_spi_com_n_247, FE_PHN293_stable_map_com_n_72, FE_PHN292_spi_com_n_43, FE_PHN291_fsm_com_n_485 : std_logic;
  signal FE_PHN290_spi_com_n_101, FE_PHN289_stable_map_com_n_98, FE_PHN288_spi_com_n_129, FE_PHN287_stable_map_com_n_111, FE_PHN286_fsm_com_n_429 : std_logic;
  signal FE_PHN285_stable_map_com_n_76, FE_PHN284_stable_map_com_n_90, FE_PHN283_stable_map_com_n_129, FE_PHN282_fsm_com_n_466, FE_PHN281_vga_com_texture_module_n_244 : std_logic;
  signal FE_PHN280_stable_map_com_n_108, FE_PHN279_spi_com_n_256, FE_PHN278_stable_map_com_n_135, FE_PHN277_stable_map_com_n_67, FE_PHN276_stable_map_com_n_71 : std_logic;
  signal FE_PHN275_spi_com_n_260, FE_PHN274_stable_map_com_n_73, FE_PHN273_stable_map_com_n_78, FE_PHN272_stable_map_com_n_56, FE_PHN271_stable_map_com_n_127 : std_logic;
  signal FE_PHN270_stable_map_com_n_68, FE_PHN269_spi_com_n_252, FE_PHN268_stable_map_com_n_128, FE_PHN267_stable_map_com_n_139, FE_PHN266_fsm_com_n_337 : std_logic;
  signal FE_PHN265_spi_com_n_175, FE_PHN264_fsm_com_n_483, FE_PHN263_stable_map_com_n_138, FE_PHN262_fsm_com_n_434, FE_PHN261_spi_com_n_182 : std_logic;
  signal FE_PHN260_spi_com_n_255, FE_PHN259_vga_com_texture_module_n_247, FE_PHN258_stable_map_com_n_92, FE_PHN257_stable_map_com_n_104, FE_PHN256_spi_com_n_261 : std_logic;
  signal FE_PHN255_spi_com_n_262, FE_PHN254_vga_com_texture_module_xposition_4, FE_PHN253_vga_com_texture_module_yposition_0, FE_PHN252_vga_com_texture_module_vvis_0, FE_PHN251_vga_com_texture_module_hvis_3 : std_logic;
  signal FE_PHN250_level_d_0, FE_PHN249_score_d_8, FE_PHN248_energy_d_4, FE_PHN247_energy_d_0, FE_PHN246_energy_d_1 : std_logic;
  signal FE_PHN245_energy_d_8, FE_PHN244_score_d_4, FE_PHN243_level_abs_0, FE_PHN242_vga_com_vcount_5, FE_PHN241_vga_com_vcount_9 : std_logic;
  signal FE_PHN240_spi_com_SCLK_count_1, FE_PHN239_vga_com_vcount_8, FE_PHN238_vga_com_vcount_7, FE_PHN237_spi_com_state_2, FE_PHN236_vga_com_hcount_8 : std_logic;
  signal FE_PHN235_vga_com_hcount_9, FE_PHN234_vga_com_vcount_6, FE_PHN233_fsm_com_n_22, FE_PHN232_energy_d_7, FE_PHN231_vga_com_vcount_2 : std_logic;
  signal FE_PHN230_fsm_com_energy_2, FE_PHN229_spi_com_SCLK_count_0, FE_PHN228_spi_com_byte_count_0, FE_PHN227_score_d_12, FE_PHN226_spi_com_bit_count_0 : std_logic;
  signal FE_PHN225_fsm_com_energy_8, FE_PHN224_fsm_com_reached_high_0, FE_PHN223_fsm_com_n_8, FE_PHN222_vga_com_display_controller_module_display_state_0, FE_PHN221_fsm_com_energy_3 : std_logic;
  signal FE_PHN220_vga_com_texture_module_n_129, FE_PHN219_vga_com_texture_module_n_134, FE_PHN218_spi_com_pause_count_0, FE_PHN217_vga_com_texture_module_n_6, FE_PHN216_vga_com_texture_module_n_115 : std_logic;
  signal FE_PHN215_fsm_com_n_6, FE_PHN214_energy_d_3, FE_PHN213_vga_com_texture_module_n_204, FE_PHN212_fsm_com_edge_detec2_3, FE_PHN211_vga_com_hcount_6 : std_logic;
  signal FE_PHN210_fsm_com_edge_detec1_3, FE_PHN209_fsm_com_edge_detec0_3, FE_PHN208_fsm_com_n_20, FE_PHN207_button_left, FE_PHN206_fsm_com_energy_7 : std_logic;
  signal FE_PHN205_fsm_com_reached_high_1, FE_PHN204_vga_com_texture_module_n_16, FE_PHN203_vga_com_texture_module_n_79, FE_PHN202_fsm_com_energy_4, FE_PHN201_n_95 : std_logic;
  signal FE_PHN200_vga_com_vcount_0, FE_PHN199_vga_com_texture_module_n_18, FE_PHN198_n_87, FE_PHN197_vga_com_texture_module_n_105, FE_PHN196_button_right : std_logic;
  signal FE_PHN195_button_up, FE_PHN194_vga_com_texture_module_n_164, FE_PHN193_vga_com_texture_module_n_17, FE_PHN192_spi_com_MOSI_shift_12, FE_PHN191_spi_com_MISO_shift_46 : std_logic;
  signal FE_PHN190_spi_com_MISO_shift_14, FE_PHN189_energy_d_2, FE_PHN188_fsm_com_n_28, FE_PHN187_spi_com_MISO_shift_12, FE_PHN186_n_93 : std_logic;
  signal FE_PHN185_spi_com_MISO_shift_34, FE_PHN184_fsm_com_n_27, FE_PHN183_map_data_volatile_33, FE_PHN182_spi_com_MOSI_shift_14, FE_PHN181_map_data_volatile_37 : std_logic;
  signal FE_PHN180_spi_com_n_5, FE_PHN179_map_data_volatile_46, FE_PHN178_map_data_volatile_36, FE_PHN177_map_data_volatile_71, FE_PHN176_stable_map_com_n_35 : std_logic;
  signal FE_PHN175_spi_com_n_9, FE_PHN174_score_d_1, FE_PHN173_spi_com_MISO_shift_11, FE_PHN172_spi_com_MISO_shift_18, FE_PHN171_map_data_10 : std_logic;
  signal FE_PHN170_spi_com_MISO_shift_40, FE_PHN169_n_86, FE_PHN168_n_91, FE_PHN167_n_94, FE_PHN166_n_90 : std_logic;
  signal FE_PHN165_n_96, FE_PHN164_n_92, FE_PHN163_n_85, FE_PHN162_spi_com_MISO_shift_3, FE_PHN161_vga_com_hcount_7 : std_logic;
  signal FE_PHN160_n_89, FE_PHN159_n_88, FE_PHN158_map_data_volatile_58, FE_PHN157_map_data_volatile_4, FE_PHN156_spi_com_MISO_shift_49 : std_logic;
  signal FE_PHN155_spi_com_MISO_shift_44, FE_PHN154_map_data_volatile_52, FE_PHN153_spi_com_MISO_shift_47, FE_PHN152_spi_com_MISO_shift_39, FE_PHN151_spi_com_MISO_shift_64 : std_logic;
  signal FE_PHN150_map_data_volatile_23, FE_PHN149_spi_com_MISO_shift_62, FE_PHN148_spi_com_MISO_shift_51, FE_PHN147_map_data_volatile_35, FE_PHN146_spi_com_MOSI_shift_5 : std_logic;
  signal FE_PHN145_spi_com_MISO_shift_27, FE_PHN144_spi_com_MISO_shift_0, FE_PHN143_fsm_com_n_12, FE_PHN142_spi_com_MOSI_shift_1, FE_PHN141_spi_com_MOSI_shift_13 : std_logic;
  signal FE_PHN140_spi_com_MISO_shift_13, FE_PHN139_map_data_volatile_53, FE_PHN138_spi_com_MISO_shift_33, FE_PHN137_map_data_volatile_16, FE_PHN136_fsm_com_edge_detec1_2 : std_logic;
  signal FE_PHN135_spi_com_MISO_shift_1, FE_PHN134_map_data_volatile_20, FE_PHN133_map_data_volatile_25, FE_PHN132_map_data_volatile_57, FE_PHN131_spi_com_MOSI_shift_7 : std_logic;
  signal FE_PHN130_map_data_volatile_38, FE_PHN129_spi_com_MOSI_shift_10, FE_PHN128_spi_com_MOSI_shift_0, FE_PHN127_map_data_volatile_3, FE_PHN126_map_data_volatile_56 : std_logic;
  signal FE_PHN125_map_data_volatile_11, FE_PHN124_map_data_volatile_8, FE_PHN123_fsm_com_edge_detec2_1, FE_PHN122_map_data_volatile_41, FE_PHN121_spi_com_MISO_shift_17 : std_logic;
  signal FE_PHN120_fsm_com_edge_detec1_1, FE_PHN119_map_data_volatile_39, FE_PHN118_map_data_volatile_45, FE_PHN117_spi_com_MISO_shift_52, FE_PHN116_map_data_volatile_9 : std_logic;
  signal FE_PHN115_spi_com_MISO_shift_61, FE_PHN114_spi_com_MISO_shift_50, FE_PHN113_map_data_volatile_62, FE_PHN112_spi_com_MOSI_shift_6, FE_PHN111_map_data_volatile_21 : std_logic;
  signal FE_PHN110_map_data_volatile_22, FE_PHN109_map_data_volatile_40, FE_PHN108_map_data_volatile_43, FE_PHN107_spi_com_MISO_shift_57, FE_PHN106_map_data_volatile_32 : std_logic;
  signal FE_PHN105_fsm_com_edge_detec0_0, FE_PHN104_map_data_volatile_61, FE_PHN103_spi_com_MISO_shift_58, FE_PHN102_spi_com_MISO_shift_65, FE_PHN101_vga_com_texture_module_vvis_6 : std_logic;
  signal FE_PHN100_fsm_com_edge_detec2_0, FE_PHN99_map_data_volatile_55, FE_PHN98_map_data_volatile_12, FE_PHN97_spi_com_MISO_shift_9, FE_PHN96_spi_com_MOSI_shift_4 : std_logic;
  signal FE_PHN95_map_data_volatile_0, FE_PHN94_map_data_volatile_6, FE_PHN93_fsm_com_edge_detec2_2, FE_PHN92_spi_com_MOSI_shift_3, FE_PHN91_fsm_com_edge_detec1_0 : std_logic;
  signal FE_PHN90_map_data_volatile_1, FE_PHN89_map_data_volatile_42, FE_PHN88_map_data_volatile_69, FE_PHN87_spi_com_MISO_shift_55, FE_PHN86_map_data_volatile_15 : std_logic;
  signal FE_PHN85_map_data_volatile_63, FE_PHN84_map_data_volatile_54, FE_PHN83_spi_com_MISO_shift_28, FE_PHN82_map_data_volatile_30, FE_PHN81_spi_com_MISO_shift_72 : std_logic;
  signal FE_PHN80_fsm_com_edge_detec0_2, FE_PHN79_fsm_com_edge_detec0_1, FE_PHN78_map_data_volatile_31, FE_PHN77_map_data_volatile_18, FE_PHN76_map_data_volatile_49 : std_logic;
  signal FE_PHN75_spi_com_MOSI_shift_2, FE_PHN74_map_data_volatile_24, FE_PHN73_map_data_volatile_47, FE_PHN72_spi_com_MISO_shift_20, FE_PHN71_map_data_volatile_5 : std_logic;
  signal FE_PHN70_map_data_volatile_66, FE_PHN69_spi_com_MISO_shift_25, FE_PHN68_spi_com_MISO_shift_10, FE_PHN67_spi_com_MISO_shift_45, FE_PHN66_spi_com_send_in0 : std_logic;
  signal FE_PHN65_map_data_volatile_50, FE_PHN64_spi_com_MISO_shift_6, FE_PHN63_map_data_volatile_26, FE_PHN62_spi_com_MISO_shift_32, FE_PHN61_map_data_volatile_17 : std_logic;
  signal FE_PHN60_map_data_volatile_67, FE_PHN59_map_data_volatile_29, FE_PHN58_map_data_volatile_70, FE_PHN57_spi_com_MISO_shift_35, FE_PHN56_map_data_volatile_34 : std_logic;
  signal FE_PHN55_map_data_volatile_14, FE_PHN54_spi_com_MISO_shift_43, FE_PHN53_spi_com_MISO_shift_26, FE_PHN52_map_data_volatile_7, FE_PHN51_spi_com_MISO_shift_41 : std_logic;
  signal FE_PHN50_map_data_volatile_48, FE_PHN49_map_data_volatile_2, FE_PHN48_map_data_volatile_68, FE_PHN47_map_data_volatile_28, FE_PHN46_spi_com_MISO_shift_4 : std_logic;
  signal FE_PHN45_map_data_volatile_59, FE_PHN44_spi_com_MISO_shift_21, FE_PHN43_map_data_volatile_19, FE_PHN42_spi_com_MISO_shift_60, FE_PHN41_map_data_volatile_27 : std_logic;
  signal FE_PHN40_spi_com_MISO_shift_29, FE_PHN39_map_data_volatile_64, FE_PHN38_map_data_volatile_60, FE_PHN37_spi_com_MISO_shift_54, FE_PHN36_map_data_volatile_13 : std_logic;
  signal FE_PHN35_spi_com_MISO_shift_22, FE_PHN34_spi_com_MISO_shift_19, FE_PHN33_map_data_volatile_65, FE_PHN32_spi_com_MISO_shift_67, FE_PHN31_spi_com_MISO_shift_48 : std_logic;
  signal FE_PHN30_spi_com_MISO_shift_15, FE_PHN29_spi_com_MISO_shift_31, FE_PHN28_spi_com_MISO_shift_68, FE_PHN27_spi_com_MISO_shift_23, FE_PHN26_spi_com_MISO_shift_59 : std_logic;
  signal FE_PHN25_spi_com_MISO_shift_38, FE_PHN24_spi_com_MISO_shift_71, FE_PHN23_spi_com_MISO_shift_24, FE_PHN22_spi_com_MISO_shift_7, FE_PHN21_spi_com_MISO_shift_70 : std_logic;
  signal FE_PHN20_spi_com_MISO_shift_36, FE_PHN19_spi_com_MISO_shift_30, FE_PHN18_spi_com_MISO_shift_2, FE_PHN17_vga_com_texture_module_n_20, FE_PHN16_spi_com_MISO_shift_66 : std_logic;
  signal FE_PHN15_spi_com_MISO_shift_53, FE_PHN14_spi_com_MISO_shift_56, FE_PHN13_spi_com_MISO_shift_69, FE_PHN12_spi_com_MISO_shift_8, FE_PHN11_spi_com_MISO_shift_37 : std_logic;
  signal FE_PHN10_spi_com_MISO_shift_16, FE_PHN9_spi_com_MISO_shift_63, FE_PHN8_spi_com_MISO_shift_5, FE_PDN7_vga_com_tile_module_n_914, FE_OFN6_spi_com_n_131 : std_logic;
  signal FE_OFN5_spi_com_n_139, FE_OFN4_vga_com_row_2, FE_OFN3_vga_com_row_1, FE_OFN2_vga_com_tile_address_0, FE_OFN1_vga_com_row_0 : std_logic;
  signal FE_OFN0_reset, CTS_24, CTS_23, CTS_22, CTS_21 : std_logic;
  signal CTS_20, CTS_19, FE_DBTN0_reset : std_logic;
  signal vga_com_display_controller_module_display_state : std_logic_vector(2 downto 0);
  signal vga_com_hcount : std_logic_vector(9 downto 0);
  signal vga_com_vcount : std_logic_vector(9 downto 0);
  signal dir_mined : std_logic_vector(2 downto 0);
  signal MOSI_data : std_logic_vector(15 downto 0);
  signal vga_com_in_red : std_logic_vector(3 downto 0);
  signal vga_com_in_blue : std_logic_vector(3 downto 0);
  signal vga_com_in_green : std_logic_vector(3 downto 0);
  signal vga_com_dim : std_logic_vector(3 downto 0);
  signal fsm_com_edge_detec2 : std_logic_vector(3 downto 0);
  signal fsm_com_edge_detec3 : std_logic_vector(3 downto 0);
  signal fsm_com_edge_detec1 : std_logic_vector(3 downto 0);
  signal map_data : std_logic_vector(71 downto 0);
  signal fsm_com_edge_detec0 : std_logic_vector(3 downto 0);
  signal game_state : std_logic_vector(1 downto 0);
  signal fsm_com_state : std_logic_vector(3 downto 0);
  signal energy_d : std_logic_vector(11 downto 0);
  signal fsm_com_energy : std_logic_vector(8 downto 0);
  signal level_d : std_logic_vector(7 downto 0);
  signal level_abs : std_logic_vector(4 downto 0);
  signal fsm_com_reached_high : std_logic_vector(1 downto 0);
  signal score_d : std_logic_vector(15 downto 0);
  signal xplayer : std_logic_vector(3 downto 0);
  signal yplayer : std_logic_vector(3 downto 0);
  signal vga_com_texture_module_vvis : std_logic_vector(6 downto 0);
  signal vga_com_texture_module_hvis : std_logic_vector(6 downto 0);
  signal vga_com_timer1 : std_logic_vector(5 downto 0);
  signal vga_com_tile_address : std_logic_vector(5 downto 0);
  signal vga_com_texture_module_frame_count : std_logic_vector(3 downto 0);
  signal vga_com_texture_module_yposition : std_logic_vector(4 downto 0);
  signal vga_com_texture_module_xposition : std_logic_vector(4 downto 0);
  signal vga_com_bg_select : std_logic_vector(2 downto 0);
  signal vga_com_column : std_logic_vector(2 downto 0);
  signal vga_com_texture_module_timer1 : std_logic_vector(5 downto 0);
  signal vga_com_row : std_logic_vector(2 downto 0);
  signal vga_com_color_address : std_logic_vector(4 downto 0);
  signal stable_map_com_state : std_logic_vector(2 downto 0);
  signal map_data_volatile : std_logic_vector(71 downto 0);
  signal spi_com_state : std_logic_vector(2 downto 0);
  signal spi_com_MISO_shift : std_logic_vector(72 downto 0);
  signal spi_com_MOSI_shift : std_logic_vector(15 downto 0);
  signal spi_com_SCLK_count : std_logic_vector(4 downto 0);
  signal spi_com_bit_count : std_logic_vector(3 downto 0);
  signal spi_com_byte_count : std_logic_vector(3 downto 0);
  signal spi_com_pause_count : std_logic_vector(2 downto 0);
  signal UNCONNECTED, UNCONNECTED0, animation_done, fsm_com_n_0, fsm_com_n_1 : std_logic;
  signal fsm_com_n_2, fsm_com_n_3, fsm_com_n_4, fsm_com_n_5, fsm_com_n_6 : std_logic;
  signal fsm_com_n_7, fsm_com_n_8, fsm_com_n_9, fsm_com_n_10, fsm_com_n_11 : std_logic;
  signal fsm_com_n_12, fsm_com_n_13, fsm_com_n_14, fsm_com_n_15, fsm_com_n_16 : std_logic;
  signal fsm_com_n_17, fsm_com_n_18, fsm_com_n_19, fsm_com_n_20, fsm_com_n_21 : std_logic;
  signal fsm_com_n_22, fsm_com_n_23, fsm_com_n_24, fsm_com_n_25, fsm_com_n_26 : std_logic;
  signal fsm_com_n_27, fsm_com_n_28, fsm_com_n_29, fsm_com_n_30, fsm_com_n_31 : std_logic;
  signal fsm_com_n_32, fsm_com_n_33, fsm_com_n_35, fsm_com_n_36, fsm_com_n_37 : std_logic;
  signal fsm_com_n_38, fsm_com_n_39, fsm_com_n_40, fsm_com_n_41, fsm_com_n_42 : std_logic;
  signal fsm_com_n_43, fsm_com_n_44, fsm_com_n_46, fsm_com_n_47, fsm_com_n_48 : std_logic;
  signal fsm_com_n_49, fsm_com_n_50, fsm_com_n_51, fsm_com_n_52, fsm_com_n_53 : std_logic;
  signal fsm_com_n_54, fsm_com_n_55, fsm_com_n_56, fsm_com_n_57, fsm_com_n_58 : std_logic;
  signal fsm_com_n_59, fsm_com_n_60, fsm_com_n_61, fsm_com_n_62, fsm_com_n_63 : std_logic;
  signal fsm_com_n_64, fsm_com_n_65, fsm_com_n_66, fsm_com_n_67, fsm_com_n_68 : std_logic;
  signal fsm_com_n_69, fsm_com_n_70, fsm_com_n_71, fsm_com_n_72, fsm_com_n_73 : std_logic;
  signal fsm_com_n_74, fsm_com_n_75, fsm_com_n_76, fsm_com_n_77, fsm_com_n_78 : std_logic;
  signal fsm_com_n_79, fsm_com_n_80, fsm_com_n_81, fsm_com_n_82, fsm_com_n_83 : std_logic;
  signal fsm_com_n_84, fsm_com_n_85, fsm_com_n_86, fsm_com_n_87, fsm_com_n_88 : std_logic;
  signal fsm_com_n_89, fsm_com_n_90, fsm_com_n_91, fsm_com_n_92, fsm_com_n_93 : std_logic;
  signal fsm_com_n_94, fsm_com_n_95, fsm_com_n_96, fsm_com_n_97, fsm_com_n_98 : std_logic;
  signal fsm_com_n_99, fsm_com_n_100, fsm_com_n_101, fsm_com_n_102, fsm_com_n_103 : std_logic;
  signal fsm_com_n_104, fsm_com_n_105, fsm_com_n_106, fsm_com_n_107, fsm_com_n_108 : std_logic;
  signal fsm_com_n_110, fsm_com_n_111, fsm_com_n_112, fsm_com_n_113, fsm_com_n_114 : std_logic;
  signal fsm_com_n_115, fsm_com_n_116, fsm_com_n_117, fsm_com_n_118, fsm_com_n_119 : std_logic;
  signal fsm_com_n_120, fsm_com_n_121, fsm_com_n_122, fsm_com_n_123, fsm_com_n_124 : std_logic;
  signal fsm_com_n_125, fsm_com_n_126, fsm_com_n_127, fsm_com_n_128, fsm_com_n_129 : std_logic;
  signal fsm_com_n_130, fsm_com_n_131, fsm_com_n_132, fsm_com_n_133, fsm_com_n_135 : std_logic;
  signal fsm_com_n_136, fsm_com_n_137, fsm_com_n_138, fsm_com_n_139, fsm_com_n_140 : std_logic;
  signal fsm_com_n_141, fsm_com_n_142, fsm_com_n_143, fsm_com_n_144, fsm_com_n_145 : std_logic;
  signal fsm_com_n_146, fsm_com_n_147, fsm_com_n_148, fsm_com_n_150, fsm_com_n_151 : std_logic;
  signal fsm_com_n_152, fsm_com_n_153, fsm_com_n_154, fsm_com_n_155, fsm_com_n_156 : std_logic;
  signal fsm_com_n_157, fsm_com_n_158, fsm_com_n_159, fsm_com_n_160, fsm_com_n_161 : std_logic;
  signal fsm_com_n_162, fsm_com_n_163, fsm_com_n_164, fsm_com_n_165, fsm_com_n_166 : std_logic;
  signal fsm_com_n_167, fsm_com_n_168, fsm_com_n_169, fsm_com_n_170, fsm_com_n_171 : std_logic;
  signal fsm_com_n_172, fsm_com_n_173, fsm_com_n_174, fsm_com_n_175, fsm_com_n_176 : std_logic;
  signal fsm_com_n_177, fsm_com_n_178, fsm_com_n_179, fsm_com_n_180, fsm_com_n_181 : std_logic;
  signal fsm_com_n_182, fsm_com_n_183, fsm_com_n_184, fsm_com_n_185, fsm_com_n_186 : std_logic;
  signal fsm_com_n_187, fsm_com_n_188, fsm_com_n_189, fsm_com_n_190, fsm_com_n_191 : std_logic;
  signal fsm_com_n_192, fsm_com_n_193, fsm_com_n_194, fsm_com_n_195, fsm_com_n_196 : std_logic;
  signal fsm_com_n_197, fsm_com_n_198, fsm_com_n_199, fsm_com_n_200, fsm_com_n_201 : std_logic;
  signal fsm_com_n_202, fsm_com_n_203, fsm_com_n_204, fsm_com_n_205, fsm_com_n_206 : std_logic;
  signal fsm_com_n_207, fsm_com_n_208, fsm_com_n_209, fsm_com_n_210, fsm_com_n_211 : std_logic;
  signal fsm_com_n_212, fsm_com_n_213, fsm_com_n_214, fsm_com_n_215, fsm_com_n_216 : std_logic;
  signal fsm_com_n_217, fsm_com_n_218, fsm_com_n_219, fsm_com_n_220, fsm_com_n_221 : std_logic;
  signal fsm_com_n_222, fsm_com_n_223, fsm_com_n_224, fsm_com_n_225, fsm_com_n_226 : std_logic;
  signal fsm_com_n_227, fsm_com_n_228, fsm_com_n_230, fsm_com_n_231, fsm_com_n_232 : std_logic;
  signal fsm_com_n_233, fsm_com_n_234, fsm_com_n_235, fsm_com_n_236, fsm_com_n_237 : std_logic;
  signal fsm_com_n_238, fsm_com_n_239, fsm_com_n_240, fsm_com_n_241, fsm_com_n_242 : std_logic;
  signal fsm_com_n_243, fsm_com_n_244, fsm_com_n_245, fsm_com_n_246, fsm_com_n_247 : std_logic;
  signal fsm_com_n_248, fsm_com_n_249, fsm_com_n_250, fsm_com_n_251, fsm_com_n_252 : std_logic;
  signal fsm_com_n_253, fsm_com_n_254, fsm_com_n_255, fsm_com_n_256, fsm_com_n_257 : std_logic;
  signal fsm_com_n_258, fsm_com_n_259, fsm_com_n_260, fsm_com_n_261, fsm_com_n_262 : std_logic;
  signal fsm_com_n_263, fsm_com_n_264, fsm_com_n_265, fsm_com_n_266, fsm_com_n_268 : std_logic;
  signal fsm_com_n_269, fsm_com_n_270, fsm_com_n_271, fsm_com_n_272, fsm_com_n_273 : std_logic;
  signal fsm_com_n_274, fsm_com_n_275, fsm_com_n_276, fsm_com_n_277, fsm_com_n_278 : std_logic;
  signal fsm_com_n_281, fsm_com_n_282, fsm_com_n_283, fsm_com_n_284, fsm_com_n_285 : std_logic;
  signal fsm_com_n_286, fsm_com_n_288, fsm_com_n_289, fsm_com_n_290, fsm_com_n_291 : std_logic;
  signal fsm_com_n_292, fsm_com_n_293, fsm_com_n_294, fsm_com_n_295, fsm_com_n_296 : std_logic;
  signal fsm_com_n_297, fsm_com_n_298, fsm_com_n_299, fsm_com_n_300, fsm_com_n_301 : std_logic;
  signal fsm_com_n_302, fsm_com_n_303, fsm_com_n_304, fsm_com_n_305, fsm_com_n_306 : std_logic;
  signal fsm_com_n_307, fsm_com_n_308, fsm_com_n_309, fsm_com_n_310, fsm_com_n_311 : std_logic;
  signal fsm_com_n_312, fsm_com_n_313, fsm_com_n_314, fsm_com_n_315, fsm_com_n_316 : std_logic;
  signal fsm_com_n_317, fsm_com_n_318, fsm_com_n_320, fsm_com_n_321, fsm_com_n_322 : std_logic;
  signal fsm_com_n_323, fsm_com_n_324, fsm_com_n_325, fsm_com_n_326, fsm_com_n_327 : std_logic;
  signal fsm_com_n_328, fsm_com_n_329, fsm_com_n_330, fsm_com_n_331, fsm_com_n_332 : std_logic;
  signal fsm_com_n_333, fsm_com_n_334, fsm_com_n_335, fsm_com_n_336, fsm_com_n_337 : std_logic;
  signal fsm_com_n_338, fsm_com_n_339, fsm_com_n_340, fsm_com_n_341, fsm_com_n_342 : std_logic;
  signal fsm_com_n_343, fsm_com_n_344, fsm_com_n_345, fsm_com_n_346, fsm_com_n_347 : std_logic;
  signal fsm_com_n_349, fsm_com_n_350, fsm_com_n_351, fsm_com_n_352, fsm_com_n_354 : std_logic;
  signal fsm_com_n_355, fsm_com_n_356, fsm_com_n_357, fsm_com_n_358, fsm_com_n_359 : std_logic;
  signal fsm_com_n_360, fsm_com_n_361, fsm_com_n_362, fsm_com_n_363, fsm_com_n_364 : std_logic;
  signal fsm_com_n_365, fsm_com_n_366, fsm_com_n_367, fsm_com_n_368, fsm_com_n_369 : std_logic;
  signal fsm_com_n_370, fsm_com_n_371, fsm_com_n_372, fsm_com_n_373, fsm_com_n_374 : std_logic;
  signal fsm_com_n_375, fsm_com_n_376, fsm_com_n_377, fsm_com_n_378, fsm_com_n_379 : std_logic;
  signal fsm_com_n_380, fsm_com_n_381, fsm_com_n_382, fsm_com_n_383, fsm_com_n_384 : std_logic;
  signal fsm_com_n_385, fsm_com_n_386, fsm_com_n_387, fsm_com_n_388, fsm_com_n_389 : std_logic;
  signal fsm_com_n_390, fsm_com_n_391, fsm_com_n_392, fsm_com_n_393, fsm_com_n_394 : std_logic;
  signal fsm_com_n_395, fsm_com_n_396, fsm_com_n_397, fsm_com_n_398, fsm_com_n_400 : std_logic;
  signal fsm_com_n_402, fsm_com_n_403, fsm_com_n_404, fsm_com_n_405, fsm_com_n_406 : std_logic;
  signal fsm_com_n_407, fsm_com_n_408, fsm_com_n_409, fsm_com_n_411, fsm_com_n_412 : std_logic;
  signal fsm_com_n_413, fsm_com_n_415, fsm_com_n_416, fsm_com_n_417, fsm_com_n_418 : std_logic;
  signal fsm_com_n_419, fsm_com_n_420, fsm_com_n_421, fsm_com_n_422, fsm_com_n_423 : std_logic;
  signal fsm_com_n_424, fsm_com_n_425, fsm_com_n_426, fsm_com_n_427, fsm_com_n_428 : std_logic;
  signal fsm_com_n_429, fsm_com_n_430, fsm_com_n_431, fsm_com_n_432, fsm_com_n_433 : std_logic;
  signal fsm_com_n_434, fsm_com_n_435, fsm_com_n_436, fsm_com_n_437, fsm_com_n_438 : std_logic;
  signal fsm_com_n_439, fsm_com_n_440, fsm_com_n_441, fsm_com_n_442, fsm_com_n_443 : std_logic;
  signal fsm_com_n_444, fsm_com_n_445, fsm_com_n_446, fsm_com_n_447, fsm_com_n_448 : std_logic;
  signal fsm_com_n_449, fsm_com_n_450, fsm_com_n_451, fsm_com_n_453, fsm_com_n_454 : std_logic;
  signal fsm_com_n_455, fsm_com_n_456, fsm_com_n_457, fsm_com_n_458, fsm_com_n_459 : std_logic;
  signal fsm_com_n_460, fsm_com_n_461, fsm_com_n_462, fsm_com_n_463, fsm_com_n_464 : std_logic;
  signal fsm_com_n_465, fsm_com_n_466, fsm_com_n_467, fsm_com_n_468, fsm_com_n_469 : std_logic;
  signal fsm_com_n_470, fsm_com_n_471, fsm_com_n_472, fsm_com_n_473, fsm_com_n_474 : std_logic;
  signal fsm_com_n_475, fsm_com_n_477, fsm_com_n_478, fsm_com_n_479, fsm_com_n_480 : std_logic;
  signal fsm_com_n_481, fsm_com_n_482, fsm_com_n_483, fsm_com_n_484, fsm_com_n_485 : std_logic;
  signal fsm_com_n_486, fsm_com_n_487, fsm_com_n_488, fsm_com_n_489, fsm_com_n_490 : std_logic;
  signal fsm_com_n_491, fsm_com_n_492, fsm_com_n_493, fsm_com_n_495, fsm_com_n_496 : std_logic;
  signal fsm_com_n_497, fsm_com_n_498, fsm_com_n_499, fsm_com_n_500, fsm_com_n_501 : std_logic;
  signal fsm_com_n_502, fsm_com_n_503, fsm_com_n_504, fsm_com_n_505, fsm_com_n_506 : std_logic;
  signal fsm_com_n_507, fsm_com_n_508, fsm_com_n_509, fsm_com_n_510, fsm_com_n_511 : std_logic;
  signal fsm_com_n_513, fsm_com_n_514, fsm_com_n_515, fsm_com_n_516, fsm_com_n_517 : std_logic;
  signal fsm_com_n_518, fsm_com_n_519, fsm_com_n_520, fsm_com_n_521, fsm_com_n_522 : std_logic;
  signal fsm_com_n_523, fsm_com_n_524, fsm_com_n_525, fsm_com_n_526, fsm_com_n_527 : std_logic;
  signal fsm_com_n_528, fsm_com_n_529, fsm_com_n_530, fsm_com_n_531, fsm_com_n_532 : std_logic;
  signal fsm_com_n_533, fsm_com_n_534, fsm_com_n_535, fsm_com_n_536, fsm_com_n_537 : std_logic;
  signal fsm_com_n_538, fsm_com_n_539, fsm_com_n_543, fsm_com_n_544, fsm_com_n_545 : std_logic;
  signal fsm_com_n_546, fsm_com_n_547, fsm_com_n_548, fsm_com_n_549, fsm_com_n_550 : std_logic;
  signal fsm_com_n_551, fsm_com_n_555, fsm_com_n_556, fsm_com_n_557, fsm_com_n_558 : std_logic;
  signal fsm_com_n_559, fsm_com_n_560, fsm_com_n_561, fsm_com_n_562, fsm_com_n_563 : std_logic;
  signal fsm_com_n_564, fsm_com_n_565, fsm_com_n_566, fsm_com_n_567, fsm_com_n_568 : std_logic;
  signal fsm_com_n_569, fsm_com_n_570, fsm_com_n_571, fsm_com_n_572, fsm_com_n_594 : std_logic;
  signal fsm_com_n_595, fsm_com_n_596, fsm_com_n_597, fsm_com_n_598, fsm_com_n_599 : std_logic;
  signal fsm_com_n_600, fsm_com_n_601, fsm_com_n_602, fsm_com_n_603, fsm_com_n_604 : std_logic;
  signal fsm_com_n_605, fsm_com_n_606, map_updated, n_0, n_1 : std_logic;
  signal n_2, n_3, n_4, n_5, n_6 : std_logic;
  signal n_7, n_8, n_9, n_10, n_11 : std_logic;
  signal n_12, n_13, n_14, n_15, n_16 : std_logic;
  signal n_17, n_18, n_19, n_20, n_21 : std_logic;
  signal n_22, n_23, n_24, n_25, n_26 : std_logic;
  signal n_27, n_28, n_29, n_30, n_31 : std_logic;
  signal n_32, n_33, n_34, n_35, n_36 : std_logic;
  signal n_37, n_38, n_39, n_40, n_41 : std_logic;
  signal n_42, n_43, n_44, n_45, n_46 : std_logic;
  signal n_47, n_48, n_49, n_50, n_51 : std_logic;
  signal n_52, n_56, n_58, n_59, n_60 : std_logic;
  signal n_61, n_62, n_63, n_64, n_65 : std_logic;
  signal n_66, n_67, n_68, n_69, n_70 : std_logic;
  signal n_71, n_72, n_73, n_74, n_75 : std_logic;
  signal n_76, n_77, n_78, n_79, n_80 : std_logic;
  signal n_81, n_82, n_83, n_84, n_85 : std_logic;
  signal n_86, n_87, n_88, n_89, n_90 : std_logic;
  signal n_91, n_92, n_93, n_94, n_95 : std_logic;
  signal n_96, n_97, n_98, n_99, n_100 : std_logic;
  signal n_101, n_102, n_103, n_104, n_105 : std_logic;
  signal n_106, n_108, n_109, n_110, n_111 : std_logic;
  signal n_112, n_116, n_142, n_143, n_144 : std_logic;
  signal n_145, n_146, send, spi_com_n_0, spi_com_n_1 : std_logic;
  signal spi_com_n_2, spi_com_n_3, spi_com_n_4, spi_com_n_5, spi_com_n_6 : std_logic;
  signal spi_com_n_7, spi_com_n_8, spi_com_n_9, spi_com_n_10, spi_com_n_12 : std_logic;
  signal spi_com_n_13, spi_com_n_14, spi_com_n_15, spi_com_n_16, spi_com_n_17 : std_logic;
  signal spi_com_n_18, spi_com_n_19, spi_com_n_20, spi_com_n_21, spi_com_n_22 : std_logic;
  signal spi_com_n_23, spi_com_n_24, spi_com_n_25, spi_com_n_26, spi_com_n_27 : std_logic;
  signal spi_com_n_28, spi_com_n_29, spi_com_n_30, spi_com_n_31, spi_com_n_32 : std_logic;
  signal spi_com_n_33, spi_com_n_34, spi_com_n_35, spi_com_n_36, spi_com_n_37 : std_logic;
  signal spi_com_n_38, spi_com_n_39, spi_com_n_40, spi_com_n_41, spi_com_n_42 : std_logic;
  signal spi_com_n_43, spi_com_n_44, spi_com_n_45, spi_com_n_46, spi_com_n_47 : std_logic;
  signal spi_com_n_48, spi_com_n_49, spi_com_n_50, spi_com_n_51, spi_com_n_52 : std_logic;
  signal spi_com_n_53, spi_com_n_54, spi_com_n_55, spi_com_n_56, spi_com_n_57 : std_logic;
  signal spi_com_n_58, spi_com_n_59, spi_com_n_60, spi_com_n_61, spi_com_n_62 : std_logic;
  signal spi_com_n_63, spi_com_n_64, spi_com_n_65, spi_com_n_66, spi_com_n_67 : std_logic;
  signal spi_com_n_68, spi_com_n_69, spi_com_n_70, spi_com_n_71, spi_com_n_72 : std_logic;
  signal spi_com_n_73, spi_com_n_74, spi_com_n_75, spi_com_n_76, spi_com_n_77 : std_logic;
  signal spi_com_n_78, spi_com_n_79, spi_com_n_80, spi_com_n_81, spi_com_n_82 : std_logic;
  signal spi_com_n_83, spi_com_n_84, spi_com_n_85, spi_com_n_86, spi_com_n_87 : std_logic;
  signal spi_com_n_88, spi_com_n_89, spi_com_n_90, spi_com_n_91, spi_com_n_92 : std_logic;
  signal spi_com_n_93, spi_com_n_94, spi_com_n_95, spi_com_n_96, spi_com_n_97 : std_logic;
  signal spi_com_n_98, spi_com_n_99, spi_com_n_100, spi_com_n_101, spi_com_n_102 : std_logic;
  signal spi_com_n_103, spi_com_n_104, spi_com_n_105, spi_com_n_106, spi_com_n_107 : std_logic;
  signal spi_com_n_108, spi_com_n_109, spi_com_n_110, spi_com_n_111, spi_com_n_112 : std_logic;
  signal spi_com_n_113, spi_com_n_114, spi_com_n_115, spi_com_n_116, spi_com_n_117 : std_logic;
  signal spi_com_n_118, spi_com_n_119, spi_com_n_120, spi_com_n_121, spi_com_n_122 : std_logic;
  signal spi_com_n_123, spi_com_n_124, spi_com_n_125, spi_com_n_126, spi_com_n_127 : std_logic;
  signal spi_com_n_128, spi_com_n_129, spi_com_n_130, spi_com_n_131, spi_com_n_132 : std_logic;
  signal spi_com_n_133, spi_com_n_134, spi_com_n_135, spi_com_n_136, spi_com_n_137 : std_logic;
  signal spi_com_n_138, spi_com_n_139, spi_com_n_140, spi_com_n_141, spi_com_n_142 : std_logic;
  signal spi_com_n_143, spi_com_n_144, spi_com_n_145, spi_com_n_146, spi_com_n_147 : std_logic;
  signal spi_com_n_148, spi_com_n_149, spi_com_n_150, spi_com_n_151, spi_com_n_152 : std_logic;
  signal spi_com_n_153, spi_com_n_154, spi_com_n_155, spi_com_n_156, spi_com_n_157 : std_logic;
  signal spi_com_n_158, spi_com_n_159, spi_com_n_160, spi_com_n_161, spi_com_n_162 : std_logic;
  signal spi_com_n_163, spi_com_n_164, spi_com_n_165, spi_com_n_166, spi_com_n_167 : std_logic;
  signal spi_com_n_168, spi_com_n_169, spi_com_n_170, spi_com_n_171, spi_com_n_172 : std_logic;
  signal spi_com_n_173, spi_com_n_174, spi_com_n_175, spi_com_n_176, spi_com_n_177 : std_logic;
  signal spi_com_n_178, spi_com_n_179, spi_com_n_180, spi_com_n_181, spi_com_n_182 : std_logic;
  signal spi_com_n_183, spi_com_n_184, spi_com_n_185, spi_com_n_186, spi_com_n_187 : std_logic;
  signal spi_com_n_188, spi_com_n_189, spi_com_n_190, spi_com_n_191, spi_com_n_192 : std_logic;
  signal spi_com_n_193, spi_com_n_194, spi_com_n_195, spi_com_n_196, spi_com_n_197 : std_logic;
  signal spi_com_n_198, spi_com_n_199, spi_com_n_200, spi_com_n_201, spi_com_n_202 : std_logic;
  signal spi_com_n_203, spi_com_n_204, spi_com_n_205, spi_com_n_206, spi_com_n_207 : std_logic;
  signal spi_com_n_208, spi_com_n_209, spi_com_n_210, spi_com_n_211, spi_com_n_212 : std_logic;
  signal spi_com_n_213, spi_com_n_214, spi_com_n_215, spi_com_n_216, spi_com_n_217 : std_logic;
  signal spi_com_n_218, spi_com_n_219, spi_com_n_220, spi_com_n_221, spi_com_n_222 : std_logic;
  signal spi_com_n_223, spi_com_n_224, spi_com_n_225, spi_com_n_226, spi_com_n_227 : std_logic;
  signal spi_com_n_228, spi_com_n_229, spi_com_n_230, spi_com_n_231, spi_com_n_232 : std_logic;
  signal spi_com_n_233, spi_com_n_234, spi_com_n_235, spi_com_n_236, spi_com_n_237 : std_logic;
  signal spi_com_n_238, spi_com_n_239, spi_com_n_240, spi_com_n_241, spi_com_n_242 : std_logic;
  signal spi_com_n_243, spi_com_n_244, spi_com_n_245, spi_com_n_246, spi_com_n_247 : std_logic;
  signal spi_com_n_248, spi_com_n_249, spi_com_n_250, spi_com_n_251, spi_com_n_252 : std_logic;
  signal spi_com_n_253, spi_com_n_254, spi_com_n_255, spi_com_n_256, spi_com_n_257 : std_logic;
  signal spi_com_n_258, spi_com_n_259, spi_com_n_260, spi_com_n_261, spi_com_n_262 : std_logic;
  signal spi_com_n_263, spi_com_n_264, spi_com_send_in0, spi_com_send_in1, stable_map_com_n_1 : std_logic;
  signal stable_map_com_n_2, stable_map_com_n_3, stable_map_com_n_4, stable_map_com_n_6, stable_map_com_n_7 : std_logic;
  signal stable_map_com_n_8, stable_map_com_n_9, stable_map_com_n_10, stable_map_com_n_11, stable_map_com_n_12 : std_logic;
  signal stable_map_com_n_13, stable_map_com_n_14, stable_map_com_n_16, stable_map_com_n_17, stable_map_com_n_18 : std_logic;
  signal stable_map_com_n_19, stable_map_com_n_20, stable_map_com_n_21, stable_map_com_n_22, stable_map_com_n_23 : std_logic;
  signal stable_map_com_n_24, stable_map_com_n_25, stable_map_com_n_26, stable_map_com_n_27, stable_map_com_n_28 : std_logic;
  signal stable_map_com_n_29, stable_map_com_n_30, stable_map_com_n_31, stable_map_com_n_32, stable_map_com_n_33 : std_logic;
  signal stable_map_com_n_34, stable_map_com_n_35, stable_map_com_n_36, stable_map_com_n_38, stable_map_com_n_39 : std_logic;
  signal stable_map_com_n_40, stable_map_com_n_41, stable_map_com_n_42, stable_map_com_n_43, stable_map_com_n_44 : std_logic;
  signal stable_map_com_n_45, stable_map_com_n_46, stable_map_com_n_47, stable_map_com_n_48, stable_map_com_n_49 : std_logic;
  signal stable_map_com_n_50, stable_map_com_n_51, stable_map_com_n_52, stable_map_com_n_53, stable_map_com_n_54 : std_logic;
  signal stable_map_com_n_55, stable_map_com_n_56, stable_map_com_n_57, stable_map_com_n_58, stable_map_com_n_59 : std_logic;
  signal stable_map_com_n_60, stable_map_com_n_61, stable_map_com_n_62, stable_map_com_n_63, stable_map_com_n_64 : std_logic;
  signal stable_map_com_n_65, stable_map_com_n_66, stable_map_com_n_67, stable_map_com_n_68, stable_map_com_n_69 : std_logic;
  signal stable_map_com_n_70, stable_map_com_n_71, stable_map_com_n_72, stable_map_com_n_73, stable_map_com_n_74 : std_logic;
  signal stable_map_com_n_75, stable_map_com_n_76, stable_map_com_n_77, stable_map_com_n_78, stable_map_com_n_79 : std_logic;
  signal stable_map_com_n_80, stable_map_com_n_81, stable_map_com_n_82, stable_map_com_n_83, stable_map_com_n_84 : std_logic;
  signal stable_map_com_n_85, stable_map_com_n_86, stable_map_com_n_87, stable_map_com_n_88, stable_map_com_n_89 : std_logic;
  signal stable_map_com_n_90, stable_map_com_n_91, stable_map_com_n_92, stable_map_com_n_93, stable_map_com_n_94 : std_logic;
  signal stable_map_com_n_95, stable_map_com_n_96, stable_map_com_n_97, stable_map_com_n_98, stable_map_com_n_99 : std_logic;
  signal stable_map_com_n_100, stable_map_com_n_101, stable_map_com_n_102, stable_map_com_n_103, stable_map_com_n_104 : std_logic;
  signal stable_map_com_n_105, stable_map_com_n_106, stable_map_com_n_107, stable_map_com_n_108, stable_map_com_n_109 : std_logic;
  signal stable_map_com_n_110, stable_map_com_n_111, stable_map_com_n_112, stable_map_com_n_113, stable_map_com_n_114 : std_logic;
  signal stable_map_com_n_115, stable_map_com_n_116, stable_map_com_n_117, stable_map_com_n_118, stable_map_com_n_119 : std_logic;
  signal stable_map_com_n_120, stable_map_com_n_121, stable_map_com_n_122, stable_map_com_n_123, stable_map_com_n_124 : std_logic;
  signal stable_map_com_n_125, stable_map_com_n_126, stable_map_com_n_127, stable_map_com_n_128, stable_map_com_n_129 : std_logic;
  signal stable_map_com_n_130, stable_map_com_n_131, stable_map_com_n_132, stable_map_com_n_133, stable_map_com_n_134 : std_logic;
  signal stable_map_com_n_135, stable_map_com_n_136, stable_map_com_n_137, stable_map_com_n_138, stable_map_com_n_139 : std_logic;
  signal stable_map_com_n_219, vga_com_color_driver_module_n_0, vga_com_color_driver_module_n_1, vga_com_color_driver_module_n_2, vga_com_color_driver_module_n_3 : std_logic;
  signal vga_com_color_driver_module_n_4, vga_com_color_driver_module_n_5, vga_com_color_driver_module_n_6, vga_com_color_driver_module_n_7, vga_com_color_driver_module_n_8 : std_logic;
  signal vga_com_color_driver_module_n_9, vga_com_color_driver_module_n_10, vga_com_color_driver_module_n_11, vga_com_color_driver_module_n_12, vga_com_color_driver_module_n_13 : std_logic;
  signal vga_com_color_driver_module_n_14, vga_com_color_driver_module_n_15, vga_com_color_driver_module_n_16, vga_com_color_driver_module_n_17, vga_com_color_driver_module_n_18 : std_logic;
  signal vga_com_color_driver_module_n_19, vga_com_color_driver_module_n_20, vga_com_color_driver_module_n_21, vga_com_color_driver_module_n_22, vga_com_color_driver_module_n_23 : std_logic;
  signal vga_com_color_driver_module_n_24, vga_com_color_driver_module_n_25, vga_com_color_driver_module_n_26, vga_com_color_driver_module_n_27, vga_com_color_driver_module_n_28 : std_logic;
  signal vga_com_color_driver_module_n_29, vga_com_color_driver_module_n_30, vga_com_color_driver_module_n_31, vga_com_color_driver_module_n_32, vga_com_color_driver_module_n_33 : std_logic;
  signal vga_com_color_driver_module_n_34, vga_com_color_driver_module_n_35, vga_com_color_driver_module_n_36, vga_com_color_driver_module_n_37, vga_com_color_driver_module_n_38 : std_logic;
  signal vga_com_color_driver_module_n_39, vga_com_color_driver_module_n_40, vga_com_color_driver_module_n_41, vga_com_color_driver_module_n_42, vga_com_color_driver_module_n_43 : std_logic;
  signal vga_com_color_driver_module_n_44, vga_com_color_driver_module_n_45, vga_com_color_driver_module_n_47, vga_com_color_driver_module_n_49, vga_com_color_driver_module_n_50 : std_logic;
  signal vga_com_color_driver_module_n_51, vga_com_color_driver_module_n_52, vga_com_color_driver_module_n_55, vga_com_texture_module_csa_tree_add_99_11_groupi_n_0, vga_com_texture_module_csa_tree_add_99_11_groupi_n_1 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_2, vga_com_texture_module_csa_tree_add_99_11_groupi_n_3, vga_com_texture_module_csa_tree_add_99_11_groupi_n_4, vga_com_texture_module_csa_tree_add_99_11_groupi_n_5, vga_com_texture_module_csa_tree_add_99_11_groupi_n_6 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_7, vga_com_texture_module_csa_tree_add_99_11_groupi_n_8, vga_com_texture_module_csa_tree_add_99_11_groupi_n_9, vga_com_texture_module_csa_tree_add_99_11_groupi_n_10, vga_com_texture_module_csa_tree_add_99_11_groupi_n_11 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_12, vga_com_texture_module_csa_tree_add_99_11_groupi_n_13, vga_com_texture_module_csa_tree_add_99_11_groupi_n_14, vga_com_texture_module_csa_tree_add_99_11_groupi_n_15, vga_com_texture_module_csa_tree_add_99_11_groupi_n_16 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_17, vga_com_texture_module_csa_tree_add_99_11_groupi_n_18, vga_com_texture_module_csa_tree_add_99_11_groupi_n_19, vga_com_texture_module_csa_tree_add_99_11_groupi_n_20, vga_com_texture_module_csa_tree_add_99_11_groupi_n_21 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_22, vga_com_texture_module_csa_tree_add_99_11_groupi_n_23, vga_com_texture_module_csa_tree_add_99_11_groupi_n_24, vga_com_texture_module_csa_tree_add_99_11_groupi_n_25, vga_com_texture_module_csa_tree_add_99_11_groupi_n_26 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_27, vga_com_texture_module_csa_tree_add_99_11_groupi_n_28, vga_com_texture_module_csa_tree_add_99_11_groupi_n_29, vga_com_texture_module_csa_tree_add_99_11_groupi_n_30, vga_com_texture_module_csa_tree_add_99_11_groupi_n_31 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_32, vga_com_texture_module_csa_tree_add_99_11_groupi_n_33, vga_com_texture_module_csa_tree_add_99_11_groupi_n_34, vga_com_texture_module_csa_tree_add_99_11_groupi_n_35, vga_com_texture_module_csa_tree_add_99_11_groupi_n_36 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_37, vga_com_texture_module_csa_tree_add_99_11_groupi_n_38, vga_com_texture_module_csa_tree_add_99_11_groupi_n_39, vga_com_texture_module_csa_tree_add_99_11_groupi_n_40, vga_com_texture_module_csa_tree_add_99_11_groupi_n_41 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_42, vga_com_texture_module_csa_tree_add_99_11_groupi_n_45, vga_com_texture_module_csa_tree_add_99_11_groupi_n_46, vga_com_texture_module_csa_tree_add_99_11_groupi_n_47, vga_com_texture_module_csa_tree_add_99_11_groupi_n_48 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_49, vga_com_texture_module_csa_tree_add_99_11_groupi_n_50, vga_com_texture_module_csa_tree_add_99_11_groupi_n_51, vga_com_texture_module_csa_tree_add_99_11_groupi_n_52, vga_com_texture_module_csa_tree_add_99_11_groupi_n_53 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_54, vga_com_texture_module_csa_tree_add_99_11_groupi_n_55, vga_com_texture_module_csa_tree_add_99_11_groupi_n_56, vga_com_texture_module_csa_tree_add_99_11_groupi_n_57, vga_com_texture_module_csa_tree_add_99_11_groupi_n_58 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_59, vga_com_texture_module_csa_tree_add_99_11_groupi_n_60, vga_com_texture_module_csa_tree_add_99_11_groupi_n_61, vga_com_texture_module_csa_tree_add_99_11_groupi_n_62, vga_com_texture_module_csa_tree_add_99_11_groupi_n_63 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_64, vga_com_texture_module_csa_tree_add_99_11_groupi_n_65, vga_com_texture_module_csa_tree_add_99_11_groupi_n_66, vga_com_texture_module_csa_tree_add_99_11_groupi_n_67, vga_com_texture_module_csa_tree_add_99_11_groupi_n_68 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_69, vga_com_texture_module_csa_tree_add_99_11_groupi_n_70, vga_com_texture_module_csa_tree_add_99_11_groupi_n_71, vga_com_texture_module_csa_tree_add_99_11_groupi_n_72, vga_com_texture_module_csa_tree_add_99_11_groupi_n_73 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_74, vga_com_texture_module_csa_tree_add_99_11_groupi_n_75, vga_com_texture_module_csa_tree_add_99_11_groupi_n_76, vga_com_texture_module_csa_tree_add_99_11_groupi_n_77, vga_com_texture_module_csa_tree_add_99_11_groupi_n_78 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_79, vga_com_texture_module_csa_tree_add_99_11_groupi_n_80, vga_com_texture_module_csa_tree_add_99_11_groupi_n_81, vga_com_texture_module_csa_tree_add_99_11_groupi_n_82, vga_com_texture_module_csa_tree_add_99_11_groupi_n_83 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_84, vga_com_texture_module_csa_tree_add_99_11_groupi_n_85, vga_com_texture_module_csa_tree_add_99_11_groupi_n_86, vga_com_texture_module_csa_tree_add_99_11_groupi_n_88, vga_com_texture_module_csa_tree_add_99_11_groupi_n_89 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_90, vga_com_texture_module_csa_tree_add_99_11_groupi_n_91, vga_com_texture_module_csa_tree_add_99_11_groupi_n_92, vga_com_texture_module_csa_tree_add_99_11_groupi_n_93, vga_com_texture_module_csa_tree_add_99_11_groupi_n_94 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_95, vga_com_texture_module_csa_tree_add_99_11_groupi_n_96, vga_com_texture_module_csa_tree_add_99_11_groupi_n_97, vga_com_texture_module_csa_tree_add_99_11_groupi_n_98, vga_com_texture_module_csa_tree_add_99_11_groupi_n_99 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_101, vga_com_texture_module_csa_tree_add_99_11_groupi_n_102, vga_com_texture_module_csa_tree_add_99_11_groupi_n_103, vga_com_texture_module_csa_tree_add_99_11_groupi_n_104, vga_com_texture_module_csa_tree_add_99_11_groupi_n_105 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_106, vga_com_texture_module_csa_tree_add_99_11_groupi_n_107, vga_com_texture_module_csa_tree_add_99_11_groupi_n_108, vga_com_texture_module_csa_tree_add_99_11_groupi_n_109, vga_com_texture_module_csa_tree_add_99_11_groupi_n_110 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_111, vga_com_texture_module_csa_tree_add_99_11_groupi_n_112, vga_com_texture_module_csa_tree_add_99_11_groupi_n_113, vga_com_texture_module_csa_tree_add_99_11_groupi_n_114, vga_com_texture_module_csa_tree_add_99_11_groupi_n_115 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_116, vga_com_texture_module_csa_tree_add_99_11_groupi_n_118, vga_com_texture_module_csa_tree_add_99_11_groupi_n_119, vga_com_texture_module_csa_tree_add_99_11_groupi_n_120, vga_com_texture_module_csa_tree_add_99_11_groupi_n_121 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_122, vga_com_texture_module_csa_tree_add_99_11_groupi_n_123, vga_com_texture_module_csa_tree_add_99_11_groupi_n_125, vga_com_texture_module_csa_tree_add_99_11_groupi_n_126, vga_com_texture_module_csa_tree_add_99_11_groupi_n_127 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_128, vga_com_texture_module_csa_tree_add_99_11_groupi_n_129, vga_com_texture_module_csa_tree_add_99_11_groupi_n_131, vga_com_texture_module_csa_tree_add_99_11_groupi_n_133, vga_com_texture_module_csa_tree_add_99_11_groupi_n_135 : std_logic;
  signal vga_com_texture_module_csa_tree_add_99_11_groupi_n_137, vga_com_texture_module_csa_tree_add_99_11_groupi_n_140, vga_com_texture_module_csa_tree_add_99_11_groupi_n_142, vga_com_texture_module_n_0, vga_com_texture_module_n_1 : std_logic;
  signal vga_com_texture_module_n_2, vga_com_texture_module_n_3, vga_com_texture_module_n_4, vga_com_texture_module_n_5, vga_com_texture_module_n_6 : std_logic;
  signal vga_com_texture_module_n_7, vga_com_texture_module_n_8, vga_com_texture_module_n_9, vga_com_texture_module_n_10, vga_com_texture_module_n_11 : std_logic;
  signal vga_com_texture_module_n_12, vga_com_texture_module_n_13, vga_com_texture_module_n_14, vga_com_texture_module_n_15, vga_com_texture_module_n_16 : std_logic;
  signal vga_com_texture_module_n_17, vga_com_texture_module_n_18, vga_com_texture_module_n_19, vga_com_texture_module_n_20, vga_com_texture_module_n_21 : std_logic;
  signal vga_com_texture_module_n_22, vga_com_texture_module_n_24, vga_com_texture_module_n_25, vga_com_texture_module_n_26, vga_com_texture_module_n_27 : std_logic;
  signal vga_com_texture_module_n_28, vga_com_texture_module_n_29, vga_com_texture_module_n_30, vga_com_texture_module_n_31, vga_com_texture_module_n_32 : std_logic;
  signal vga_com_texture_module_n_33, vga_com_texture_module_n_34, vga_com_texture_module_n_35, vga_com_texture_module_n_36, vga_com_texture_module_n_37 : std_logic;
  signal vga_com_texture_module_n_38, vga_com_texture_module_n_39, vga_com_texture_module_n_40, vga_com_texture_module_n_41, vga_com_texture_module_n_42 : std_logic;
  signal vga_com_texture_module_n_43, vga_com_texture_module_n_44, vga_com_texture_module_n_45, vga_com_texture_module_n_46, vga_com_texture_module_n_47 : std_logic;
  signal vga_com_texture_module_n_48, vga_com_texture_module_n_49, vga_com_texture_module_n_50, vga_com_texture_module_n_51, vga_com_texture_module_n_52 : std_logic;
  signal vga_com_texture_module_n_53, vga_com_texture_module_n_54, vga_com_texture_module_n_55, vga_com_texture_module_n_56, vga_com_texture_module_n_57 : std_logic;
  signal vga_com_texture_module_n_58, vga_com_texture_module_n_59, vga_com_texture_module_n_60, vga_com_texture_module_n_61, vga_com_texture_module_n_62 : std_logic;
  signal vga_com_texture_module_n_63, vga_com_texture_module_n_64, vga_com_texture_module_n_65, vga_com_texture_module_n_66, vga_com_texture_module_n_67 : std_logic;
  signal vga_com_texture_module_n_68, vga_com_texture_module_n_69, vga_com_texture_module_n_70, vga_com_texture_module_n_71, vga_com_texture_module_n_72 : std_logic;
  signal vga_com_texture_module_n_73, vga_com_texture_module_n_74, vga_com_texture_module_n_75, vga_com_texture_module_n_76, vga_com_texture_module_n_77 : std_logic;
  signal vga_com_texture_module_n_78, vga_com_texture_module_n_79, vga_com_texture_module_n_80, vga_com_texture_module_n_81, vga_com_texture_module_n_82 : std_logic;
  signal vga_com_texture_module_n_83, vga_com_texture_module_n_84, vga_com_texture_module_n_85, vga_com_texture_module_n_86, vga_com_texture_module_n_87 : std_logic;
  signal vga_com_texture_module_n_88, vga_com_texture_module_n_89, vga_com_texture_module_n_90, vga_com_texture_module_n_91, vga_com_texture_module_n_92 : std_logic;
  signal vga_com_texture_module_n_93, vga_com_texture_module_n_94, vga_com_texture_module_n_95, vga_com_texture_module_n_96, vga_com_texture_module_n_97 : std_logic;
  signal vga_com_texture_module_n_98, vga_com_texture_module_n_99, vga_com_texture_module_n_100, vga_com_texture_module_n_101, vga_com_texture_module_n_102 : std_logic;
  signal vga_com_texture_module_n_103, vga_com_texture_module_n_104, vga_com_texture_module_n_105, vga_com_texture_module_n_106, vga_com_texture_module_n_107 : std_logic;
  signal vga_com_texture_module_n_108, vga_com_texture_module_n_109, vga_com_texture_module_n_110, vga_com_texture_module_n_111, vga_com_texture_module_n_112 : std_logic;
  signal vga_com_texture_module_n_113, vga_com_texture_module_n_114, vga_com_texture_module_n_115, vga_com_texture_module_n_116, vga_com_texture_module_n_117 : std_logic;
  signal vga_com_texture_module_n_118, vga_com_texture_module_n_119, vga_com_texture_module_n_120, vga_com_texture_module_n_121, vga_com_texture_module_n_122 : std_logic;
  signal vga_com_texture_module_n_123, vga_com_texture_module_n_124, vga_com_texture_module_n_125, vga_com_texture_module_n_126, vga_com_texture_module_n_127 : std_logic;
  signal vga_com_texture_module_n_128, vga_com_texture_module_n_129, vga_com_texture_module_n_130, vga_com_texture_module_n_131, vga_com_texture_module_n_132 : std_logic;
  signal vga_com_texture_module_n_133, vga_com_texture_module_n_134, vga_com_texture_module_n_135, vga_com_texture_module_n_136, vga_com_texture_module_n_137 : std_logic;
  signal vga_com_texture_module_n_138, vga_com_texture_module_n_139, vga_com_texture_module_n_140, vga_com_texture_module_n_141, vga_com_texture_module_n_142 : std_logic;
  signal vga_com_texture_module_n_143, vga_com_texture_module_n_144, vga_com_texture_module_n_145, vga_com_texture_module_n_146, vga_com_texture_module_n_147 : std_logic;
  signal vga_com_texture_module_n_148, vga_com_texture_module_n_149, vga_com_texture_module_n_150, vga_com_texture_module_n_151, vga_com_texture_module_n_152 : std_logic;
  signal vga_com_texture_module_n_153, vga_com_texture_module_n_154, vga_com_texture_module_n_155, vga_com_texture_module_n_156, vga_com_texture_module_n_157 : std_logic;
  signal vga_com_texture_module_n_158, vga_com_texture_module_n_159, vga_com_texture_module_n_160, vga_com_texture_module_n_161, vga_com_texture_module_n_162 : std_logic;
  signal vga_com_texture_module_n_163, vga_com_texture_module_n_164, vga_com_texture_module_n_165, vga_com_texture_module_n_166, vga_com_texture_module_n_167 : std_logic;
  signal vga_com_texture_module_n_168, vga_com_texture_module_n_169, vga_com_texture_module_n_170, vga_com_texture_module_n_171, vga_com_texture_module_n_172 : std_logic;
  signal vga_com_texture_module_n_173, vga_com_texture_module_n_174, vga_com_texture_module_n_175, vga_com_texture_module_n_176, vga_com_texture_module_n_177 : std_logic;
  signal vga_com_texture_module_n_178, vga_com_texture_module_n_179, vga_com_texture_module_n_180, vga_com_texture_module_n_181, vga_com_texture_module_n_182 : std_logic;
  signal vga_com_texture_module_n_183, vga_com_texture_module_n_184, vga_com_texture_module_n_185, vga_com_texture_module_n_186, vga_com_texture_module_n_187 : std_logic;
  signal vga_com_texture_module_n_188, vga_com_texture_module_n_189, vga_com_texture_module_n_190, vga_com_texture_module_n_191, vga_com_texture_module_n_192 : std_logic;
  signal vga_com_texture_module_n_193, vga_com_texture_module_n_194, vga_com_texture_module_n_195, vga_com_texture_module_n_196, vga_com_texture_module_n_197 : std_logic;
  signal vga_com_texture_module_n_198, vga_com_texture_module_n_199, vga_com_texture_module_n_200, vga_com_texture_module_n_201, vga_com_texture_module_n_202 : std_logic;
  signal vga_com_texture_module_n_203, vga_com_texture_module_n_204, vga_com_texture_module_n_205, vga_com_texture_module_n_206, vga_com_texture_module_n_207 : std_logic;
  signal vga_com_texture_module_n_208, vga_com_texture_module_n_209, vga_com_texture_module_n_210, vga_com_texture_module_n_211, vga_com_texture_module_n_212 : std_logic;
  signal vga_com_texture_module_n_213, vga_com_texture_module_n_214, vga_com_texture_module_n_215, vga_com_texture_module_n_216, vga_com_texture_module_n_217 : std_logic;
  signal vga_com_texture_module_n_218, vga_com_texture_module_n_219, vga_com_texture_module_n_220, vga_com_texture_module_n_221, vga_com_texture_module_n_222 : std_logic;
  signal vga_com_texture_module_n_223, vga_com_texture_module_n_224, vga_com_texture_module_n_225, vga_com_texture_module_n_226, vga_com_texture_module_n_227 : std_logic;
  signal vga_com_texture_module_n_228, vga_com_texture_module_n_229, vga_com_texture_module_n_230, vga_com_texture_module_n_231, vga_com_texture_module_n_232 : std_logic;
  signal vga_com_texture_module_n_233, vga_com_texture_module_n_234, vga_com_texture_module_n_235, vga_com_texture_module_n_236, vga_com_texture_module_n_237 : std_logic;
  signal vga_com_texture_module_n_238, vga_com_texture_module_n_239, vga_com_texture_module_n_240, vga_com_texture_module_n_241, vga_com_texture_module_n_242 : std_logic;
  signal vga_com_texture_module_n_243, vga_com_texture_module_n_244, vga_com_texture_module_n_245, vga_com_texture_module_n_246, vga_com_texture_module_n_247 : std_logic;
  signal vga_com_texture_module_n_248, vga_com_texture_module_n_249, vga_com_texture_module_n_250, vga_com_texture_module_n_251, vga_com_texture_module_n_252 : std_logic;
  signal vga_com_texture_module_n_253, vga_com_texture_module_n_254, vga_com_texture_module_n_256, vga_com_texture_module_n_257, vga_com_texture_module_n_259 : std_logic;
  signal vga_com_texture_module_n_260, vga_com_texture_module_n_262, vga_com_texture_module_n_263, vga_com_texture_module_n_264, vga_com_texture_module_n_265 : std_logic;
  signal vga_com_texture_module_n_266, vga_com_texture_module_n_267, vga_com_texture_module_n_268, vga_com_texture_module_n_269, vga_com_texture_module_n_270 : std_logic;
  signal vga_com_texture_module_n_271, vga_com_texture_module_n_272, vga_com_texture_module_n_273, vga_com_texture_module_n_274, vga_com_texture_module_n_275 : std_logic;
  signal vga_com_texture_module_n_276, vga_com_texture_module_n_277, vga_com_texture_module_n_278, vga_com_texture_module_n_279, vga_com_texture_module_n_280 : std_logic;
  signal vga_com_texture_module_n_281, vga_com_texture_module_n_282, vga_com_texture_module_n_283, vga_com_texture_module_n_285, vga_com_texture_module_n_286 : std_logic;
  signal vga_com_texture_module_n_287, vga_com_texture_module_n_288, vga_com_texture_module_n_289, vga_com_texture_module_n_290, vga_com_texture_module_n_291 : std_logic;
  signal vga_com_texture_module_n_292, vga_com_texture_module_n_293, vga_com_texture_module_n_294, vga_com_texture_module_n_295, vga_com_texture_module_n_296 : std_logic;
  signal vga_com_texture_module_n_297, vga_com_texture_module_n_298, vga_com_texture_module_n_299, vga_com_texture_module_n_300, vga_com_texture_module_n_301 : std_logic;
  signal vga_com_texture_module_n_302, vga_com_texture_module_n_303, vga_com_texture_module_n_304, vga_com_texture_module_n_305, vga_com_texture_module_n_306 : std_logic;
  signal vga_com_texture_module_n_307, vga_com_texture_module_n_308, vga_com_texture_module_n_309, vga_com_texture_module_n_310, vga_com_texture_module_n_311 : std_logic;
  signal vga_com_texture_module_n_312, vga_com_texture_module_n_313, vga_com_texture_module_n_314, vga_com_texture_module_n_315, vga_com_texture_module_n_316 : std_logic;
  signal vga_com_texture_module_n_317, vga_com_texture_module_n_318, vga_com_texture_module_n_319, vga_com_texture_module_n_320, vga_com_texture_module_n_321 : std_logic;
  signal vga_com_texture_module_n_322, vga_com_texture_module_n_323, vga_com_texture_module_n_324, vga_com_texture_module_n_325, vga_com_texture_module_n_326 : std_logic;
  signal vga_com_texture_module_n_327, vga_com_texture_module_n_328, vga_com_texture_module_n_329, vga_com_texture_module_n_330, vga_com_texture_module_n_331 : std_logic;
  signal vga_com_texture_module_n_332, vga_com_texture_module_n_333, vga_com_texture_module_n_334, vga_com_texture_module_n_335, vga_com_texture_module_n_336 : std_logic;
  signal vga_com_texture_module_n_337, vga_com_texture_module_n_338, vga_com_texture_module_n_339, vga_com_texture_module_n_340, vga_com_texture_module_n_341 : std_logic;
  signal vga_com_texture_module_n_342, vga_com_texture_module_n_343, vga_com_texture_module_n_344, vga_com_texture_module_n_345, vga_com_texture_module_n_346 : std_logic;
  signal vga_com_texture_module_n_347, vga_com_texture_module_n_348, vga_com_texture_module_n_349, vga_com_texture_module_n_350, vga_com_texture_module_n_351 : std_logic;
  signal vga_com_texture_module_n_352, vga_com_texture_module_n_353, vga_com_texture_module_n_354, vga_com_texture_module_n_355, vga_com_texture_module_n_356 : std_logic;
  signal vga_com_texture_module_n_357, vga_com_texture_module_n_358, vga_com_texture_module_n_359, vga_com_texture_module_n_360, vga_com_texture_module_n_361 : std_logic;
  signal vga_com_texture_module_n_362, vga_com_texture_module_n_363, vga_com_texture_module_n_364, vga_com_texture_module_n_365, vga_com_texture_module_n_366 : std_logic;
  signal vga_com_texture_module_n_367, vga_com_texture_module_n_368, vga_com_texture_module_n_369, vga_com_texture_module_n_370, vga_com_texture_module_n_371 : std_logic;
  signal vga_com_texture_module_n_372, vga_com_texture_module_n_373, vga_com_texture_module_n_374, vga_com_texture_module_n_375, vga_com_texture_module_n_376 : std_logic;
  signal vga_com_texture_module_n_377, vga_com_texture_module_n_378, vga_com_texture_module_n_379, vga_com_texture_module_n_380, vga_com_texture_module_n_381 : std_logic;
  signal vga_com_texture_module_n_382, vga_com_texture_module_n_383, vga_com_texture_module_n_384, vga_com_texture_module_n_385, vga_com_texture_module_n_386 : std_logic;
  signal vga_com_texture_module_n_387, vga_com_texture_module_n_388, vga_com_texture_module_n_389, vga_com_texture_module_n_390, vga_com_texture_module_n_391 : std_logic;
  signal vga_com_texture_module_n_392, vga_com_texture_module_n_393, vga_com_texture_module_n_394, vga_com_texture_module_n_395, vga_com_texture_module_n_396 : std_logic;
  signal vga_com_texture_module_n_397, vga_com_texture_module_n_398, vga_com_texture_module_n_399, vga_com_texture_module_n_400, vga_com_texture_module_n_401 : std_logic;
  signal vga_com_texture_module_n_402, vga_com_texture_module_n_403, vga_com_texture_module_n_404, vga_com_texture_module_n_405, vga_com_texture_module_n_406 : std_logic;
  signal vga_com_texture_module_n_407, vga_com_texture_module_n_408, vga_com_texture_module_n_409, vga_com_texture_module_n_410, vga_com_texture_module_n_411 : std_logic;
  signal vga_com_texture_module_n_412, vga_com_texture_module_n_413, vga_com_texture_module_n_414, vga_com_texture_module_n_415, vga_com_texture_module_n_416 : std_logic;
  signal vga_com_texture_module_n_417, vga_com_texture_module_n_418, vga_com_texture_module_n_419, vga_com_texture_module_n_420, vga_com_texture_module_n_421 : std_logic;
  signal vga_com_texture_module_n_422, vga_com_texture_module_n_423, vga_com_texture_module_n_424, vga_com_texture_module_n_425, vga_com_texture_module_n_426 : std_logic;
  signal vga_com_texture_module_n_427, vga_com_texture_module_n_428, vga_com_texture_module_n_429, vga_com_texture_module_n_430, vga_com_texture_module_n_431 : std_logic;
  signal vga_com_texture_module_n_432, vga_com_texture_module_n_433, vga_com_texture_module_n_434, vga_com_texture_module_n_435, vga_com_texture_module_n_436 : std_logic;
  signal vga_com_texture_module_n_437, vga_com_texture_module_n_438, vga_com_texture_module_n_439, vga_com_texture_module_n_440, vga_com_texture_module_n_441 : std_logic;
  signal vga_com_texture_module_n_442, vga_com_texture_module_n_443, vga_com_texture_module_n_444, vga_com_texture_module_n_445, vga_com_texture_module_n_446 : std_logic;
  signal vga_com_texture_module_n_447, vga_com_texture_module_n_448, vga_com_texture_module_n_449, vga_com_texture_module_n_450, vga_com_texture_module_n_451 : std_logic;
  signal vga_com_texture_module_n_452, vga_com_texture_module_n_453, vga_com_texture_module_n_454, vga_com_texture_module_n_455, vga_com_texture_module_n_456 : std_logic;
  signal vga_com_texture_module_n_457, vga_com_texture_module_n_458, vga_com_texture_module_n_459, vga_com_texture_module_n_460, vga_com_texture_module_n_461 : std_logic;
  signal vga_com_texture_module_n_462, vga_com_texture_module_n_463, vga_com_texture_module_n_464, vga_com_texture_module_n_465, vga_com_texture_module_n_466 : std_logic;
  signal vga_com_texture_module_n_467, vga_com_texture_module_n_468, vga_com_texture_module_n_469, vga_com_texture_module_n_470, vga_com_texture_module_n_471 : std_logic;
  signal vga_com_texture_module_n_472, vga_com_texture_module_n_473, vga_com_texture_module_n_474, vga_com_texture_module_n_475, vga_com_texture_module_n_476 : std_logic;
  signal vga_com_texture_module_n_477, vga_com_texture_module_n_478, vga_com_texture_module_n_479, vga_com_texture_module_n_480, vga_com_texture_module_n_481 : std_logic;
  signal vga_com_texture_module_n_482, vga_com_texture_module_n_483, vga_com_texture_module_n_484, vga_com_texture_module_n_485, vga_com_texture_module_n_486 : std_logic;
  signal vga_com_texture_module_n_487, vga_com_texture_module_n_488, vga_com_texture_module_n_489, vga_com_texture_module_n_490, vga_com_texture_module_n_491 : std_logic;
  signal vga_com_texture_module_n_492, vga_com_texture_module_n_493, vga_com_texture_module_n_494, vga_com_texture_module_n_495, vga_com_texture_module_n_496 : std_logic;
  signal vga_com_texture_module_n_497, vga_com_texture_module_n_498, vga_com_texture_module_n_499, vga_com_texture_module_n_500, vga_com_texture_module_n_501 : std_logic;
  signal vga_com_texture_module_n_502, vga_com_texture_module_n_503, vga_com_texture_module_n_504, vga_com_texture_module_n_505, vga_com_texture_module_n_506 : std_logic;
  signal vga_com_texture_module_n_507, vga_com_texture_module_n_508, vga_com_texture_module_n_509, vga_com_texture_module_n_510, vga_com_texture_module_n_511 : std_logic;
  signal vga_com_texture_module_n_512, vga_com_texture_module_n_513, vga_com_texture_module_n_514, vga_com_texture_module_n_515, vga_com_texture_module_n_516 : std_logic;
  signal vga_com_texture_module_n_517, vga_com_texture_module_n_518, vga_com_texture_module_n_519, vga_com_texture_module_n_520, vga_com_texture_module_n_521 : std_logic;
  signal vga_com_texture_module_n_522, vga_com_texture_module_n_523, vga_com_texture_module_n_524, vga_com_texture_module_n_525, vga_com_texture_module_n_526 : std_logic;
  signal vga_com_texture_module_n_527, vga_com_texture_module_n_528, vga_com_texture_module_n_529, vga_com_texture_module_n_530, vga_com_texture_module_n_531 : std_logic;
  signal vga_com_texture_module_n_532, vga_com_texture_module_n_533, vga_com_texture_module_n_534, vga_com_texture_module_n_535, vga_com_texture_module_n_536 : std_logic;
  signal vga_com_texture_module_n_537, vga_com_texture_module_n_538, vga_com_texture_module_n_539, vga_com_texture_module_n_540, vga_com_texture_module_n_541 : std_logic;
  signal vga_com_texture_module_n_542, vga_com_texture_module_n_543, vga_com_texture_module_n_544, vga_com_texture_module_n_545, vga_com_texture_module_n_546 : std_logic;
  signal vga_com_texture_module_n_547, vga_com_texture_module_n_548, vga_com_texture_module_n_549, vga_com_texture_module_n_550, vga_com_texture_module_n_551 : std_logic;
  signal vga_com_texture_module_n_552, vga_com_texture_module_n_553, vga_com_texture_module_n_554, vga_com_texture_module_n_555, vga_com_texture_module_n_556 : std_logic;
  signal vga_com_texture_module_n_557, vga_com_texture_module_n_558, vga_com_texture_module_n_559, vga_com_texture_module_n_560, vga_com_texture_module_n_561 : std_logic;
  signal vga_com_texture_module_n_562, vga_com_texture_module_n_563, vga_com_texture_module_n_564, vga_com_texture_module_n_565, vga_com_texture_module_n_566 : std_logic;
  signal vga_com_texture_module_n_567, vga_com_texture_module_n_568, vga_com_texture_module_n_569, vga_com_texture_module_n_570, vga_com_texture_module_n_571 : std_logic;
  signal vga_com_texture_module_n_572, vga_com_texture_module_n_573, vga_com_texture_module_n_574, vga_com_texture_module_n_575, vga_com_texture_module_n_576 : std_logic;
  signal vga_com_texture_module_n_577, vga_com_texture_module_n_578, vga_com_texture_module_n_579, vga_com_texture_module_n_580, vga_com_texture_module_n_581 : std_logic;
  signal vga_com_texture_module_n_582, vga_com_texture_module_n_583, vga_com_texture_module_n_584, vga_com_texture_module_n_585, vga_com_texture_module_n_586 : std_logic;
  signal vga_com_texture_module_n_587, vga_com_texture_module_n_588, vga_com_texture_module_n_589, vga_com_texture_module_n_590, vga_com_texture_module_n_591 : std_logic;
  signal vga_com_texture_module_n_592, vga_com_texture_module_n_593, vga_com_texture_module_n_594, vga_com_texture_module_n_595, vga_com_texture_module_n_596 : std_logic;
  signal vga_com_texture_module_n_597, vga_com_texture_module_n_598, vga_com_texture_module_n_599, vga_com_texture_module_n_600, vga_com_texture_module_n_601 : std_logic;
  signal vga_com_texture_module_n_602, vga_com_texture_module_n_603, vga_com_texture_module_n_604, vga_com_texture_module_n_605, vga_com_texture_module_n_606 : std_logic;
  signal vga_com_texture_module_n_607, vga_com_texture_module_n_608, vga_com_texture_module_n_609, vga_com_texture_module_n_610, vga_com_texture_module_n_611 : std_logic;
  signal vga_com_texture_module_n_612, vga_com_texture_module_n_613, vga_com_texture_module_n_614, vga_com_texture_module_n_615, vga_com_texture_module_n_616 : std_logic;
  signal vga_com_texture_module_n_617, vga_com_texture_module_n_618, vga_com_texture_module_n_619, vga_com_texture_module_n_620, vga_com_texture_module_n_621 : std_logic;
  signal vga_com_texture_module_n_622, vga_com_texture_module_n_623, vga_com_texture_module_n_624, vga_com_texture_module_n_625, vga_com_texture_module_n_626 : std_logic;
  signal vga_com_texture_module_n_627, vga_com_texture_module_n_628, vga_com_texture_module_n_629, vga_com_texture_module_n_630, vga_com_texture_module_n_631 : std_logic;
  signal vga_com_texture_module_n_632, vga_com_texture_module_n_633, vga_com_texture_module_n_634, vga_com_texture_module_n_635, vga_com_texture_module_n_636 : std_logic;
  signal vga_com_texture_module_n_637, vga_com_texture_module_n_638, vga_com_texture_module_n_639, vga_com_texture_module_n_640, vga_com_texture_module_n_641 : std_logic;
  signal vga_com_texture_module_n_642, vga_com_texture_module_n_643, vga_com_texture_module_n_644, vga_com_texture_module_n_645, vga_com_texture_module_n_646 : std_logic;
  signal vga_com_texture_module_n_647, vga_com_texture_module_n_648, vga_com_texture_module_n_650, vga_com_texture_module_n_651, vga_com_texture_module_n_652 : std_logic;
  signal vga_com_texture_module_n_653, vga_com_texture_module_n_654, vga_com_texture_module_n_655, vga_com_texture_module_n_656, vga_com_texture_module_n_657 : std_logic;
  signal vga_com_texture_module_n_658, vga_com_texture_module_n_659, vga_com_texture_module_n_660, vga_com_texture_module_n_661, vga_com_texture_module_n_662 : std_logic;
  signal vga_com_texture_module_n_663, vga_com_texture_module_n_664, vga_com_texture_module_n_667, vga_com_texture_module_n_668, vga_com_texture_module_n_669 : std_logic;
  signal vga_com_texture_module_n_670, vga_com_texture_module_n_671, vga_com_texture_module_n_672, vga_com_texture_module_n_673, vga_com_texture_module_n_674 : std_logic;
  signal vga_com_texture_module_n_675, vga_com_texture_module_n_676, vga_com_texture_module_n_678, vga_com_texture_module_n_679, vga_com_texture_module_n_681 : std_logic;
  signal vga_com_texture_module_n_682, vga_com_texture_module_n_683, vga_com_texture_module_n_684, vga_com_texture_module_n_685, vga_com_texture_module_n_686 : std_logic;
  signal vga_com_texture_module_n_687, vga_com_texture_module_n_688, vga_com_texture_module_n_689, vga_com_texture_module_n_690, vga_com_texture_module_n_691 : std_logic;
  signal vga_com_texture_module_n_692, vga_com_texture_module_n_693, vga_com_texture_module_n_694, vga_com_texture_module_n_695, vga_com_texture_module_n_696 : std_logic;
  signal vga_com_texture_module_n_697, vga_com_texture_module_n_698, vga_com_texture_module_n_699, vga_com_texture_module_n_700, vga_com_texture_module_n_701 : std_logic;
  signal vga_com_texture_module_n_702, vga_com_texture_module_n_703, vga_com_texture_module_n_705, vga_com_texture_module_n_706, vga_com_texture_module_n_707 : std_logic;
  signal vga_com_texture_module_n_708, vga_com_texture_module_n_709, vga_com_texture_module_n_710, vga_com_texture_module_n_711, vga_com_texture_module_n_712 : std_logic;
  signal vga_com_texture_module_n_850, vga_com_tile_module_n_0, vga_com_tile_module_n_1, vga_com_tile_module_n_2, vga_com_tile_module_n_3 : std_logic;
  signal vga_com_tile_module_n_4, vga_com_tile_module_n_5, vga_com_tile_module_n_6, vga_com_tile_module_n_7, vga_com_tile_module_n_8 : std_logic;
  signal vga_com_tile_module_n_9, vga_com_tile_module_n_10, vga_com_tile_module_n_11, vga_com_tile_module_n_12, vga_com_tile_module_n_13 : std_logic;
  signal vga_com_tile_module_n_14, vga_com_tile_module_n_15, vga_com_tile_module_n_16, vga_com_tile_module_n_17, vga_com_tile_module_n_18 : std_logic;
  signal vga_com_tile_module_n_19, vga_com_tile_module_n_20, vga_com_tile_module_n_21, vga_com_tile_module_n_22, vga_com_tile_module_n_23 : std_logic;
  signal vga_com_tile_module_n_24, vga_com_tile_module_n_25, vga_com_tile_module_n_26, vga_com_tile_module_n_27, vga_com_tile_module_n_28 : std_logic;
  signal vga_com_tile_module_n_29, vga_com_tile_module_n_30, vga_com_tile_module_n_31, vga_com_tile_module_n_32, vga_com_tile_module_n_33 : std_logic;
  signal vga_com_tile_module_n_34, vga_com_tile_module_n_35, vga_com_tile_module_n_36, vga_com_tile_module_n_37, vga_com_tile_module_n_38 : std_logic;
  signal vga_com_tile_module_n_39, vga_com_tile_module_n_40, vga_com_tile_module_n_41, vga_com_tile_module_n_42, vga_com_tile_module_n_43 : std_logic;
  signal vga_com_tile_module_n_44, vga_com_tile_module_n_45, vga_com_tile_module_n_46, vga_com_tile_module_n_47, vga_com_tile_module_n_48 : std_logic;
  signal vga_com_tile_module_n_49, vga_com_tile_module_n_50, vga_com_tile_module_n_51, vga_com_tile_module_n_52, vga_com_tile_module_n_53 : std_logic;
  signal vga_com_tile_module_n_54, vga_com_tile_module_n_55, vga_com_tile_module_n_56, vga_com_tile_module_n_57, vga_com_tile_module_n_58 : std_logic;
  signal vga_com_tile_module_n_59, vga_com_tile_module_n_60, vga_com_tile_module_n_61, vga_com_tile_module_n_62, vga_com_tile_module_n_63 : std_logic;
  signal vga_com_tile_module_n_64, vga_com_tile_module_n_65, vga_com_tile_module_n_66, vga_com_tile_module_n_67, vga_com_tile_module_n_68 : std_logic;
  signal vga_com_tile_module_n_69, vga_com_tile_module_n_70, vga_com_tile_module_n_71, vga_com_tile_module_n_72, vga_com_tile_module_n_73 : std_logic;
  signal vga_com_tile_module_n_74, vga_com_tile_module_n_75, vga_com_tile_module_n_76, vga_com_tile_module_n_77, vga_com_tile_module_n_78 : std_logic;
  signal vga_com_tile_module_n_79, vga_com_tile_module_n_80, vga_com_tile_module_n_81, vga_com_tile_module_n_82, vga_com_tile_module_n_83 : std_logic;
  signal vga_com_tile_module_n_84, vga_com_tile_module_n_85, vga_com_tile_module_n_86, vga_com_tile_module_n_87, vga_com_tile_module_n_88 : std_logic;
  signal vga_com_tile_module_n_89, vga_com_tile_module_n_90, vga_com_tile_module_n_91, vga_com_tile_module_n_92, vga_com_tile_module_n_93 : std_logic;
  signal vga_com_tile_module_n_94, vga_com_tile_module_n_95, vga_com_tile_module_n_96, vga_com_tile_module_n_97, vga_com_tile_module_n_98 : std_logic;
  signal vga_com_tile_module_n_99, vga_com_tile_module_n_100, vga_com_tile_module_n_101, vga_com_tile_module_n_102, vga_com_tile_module_n_103 : std_logic;
  signal vga_com_tile_module_n_104, vga_com_tile_module_n_105, vga_com_tile_module_n_106, vga_com_tile_module_n_107, vga_com_tile_module_n_108 : std_logic;
  signal vga_com_tile_module_n_109, vga_com_tile_module_n_110, vga_com_tile_module_n_111, vga_com_tile_module_n_112, vga_com_tile_module_n_113 : std_logic;
  signal vga_com_tile_module_n_114, vga_com_tile_module_n_115, vga_com_tile_module_n_116, vga_com_tile_module_n_117, vga_com_tile_module_n_118 : std_logic;
  signal vga_com_tile_module_n_119, vga_com_tile_module_n_120, vga_com_tile_module_n_121, vga_com_tile_module_n_122, vga_com_tile_module_n_123 : std_logic;
  signal vga_com_tile_module_n_124, vga_com_tile_module_n_125, vga_com_tile_module_n_126, vga_com_tile_module_n_127, vga_com_tile_module_n_128 : std_logic;
  signal vga_com_tile_module_n_129, vga_com_tile_module_n_130, vga_com_tile_module_n_131, vga_com_tile_module_n_132, vga_com_tile_module_n_133 : std_logic;
  signal vga_com_tile_module_n_134, vga_com_tile_module_n_135, vga_com_tile_module_n_136, vga_com_tile_module_n_137, vga_com_tile_module_n_138 : std_logic;
  signal vga_com_tile_module_n_139, vga_com_tile_module_n_140, vga_com_tile_module_n_141, vga_com_tile_module_n_142, vga_com_tile_module_n_143 : std_logic;
  signal vga_com_tile_module_n_144, vga_com_tile_module_n_145, vga_com_tile_module_n_146, vga_com_tile_module_n_147, vga_com_tile_module_n_148 : std_logic;
  signal vga_com_tile_module_n_149, vga_com_tile_module_n_150, vga_com_tile_module_n_151, vga_com_tile_module_n_152, vga_com_tile_module_n_153 : std_logic;
  signal vga_com_tile_module_n_154, vga_com_tile_module_n_155, vga_com_tile_module_n_156, vga_com_tile_module_n_157, vga_com_tile_module_n_158 : std_logic;
  signal vga_com_tile_module_n_159, vga_com_tile_module_n_160, vga_com_tile_module_n_161, vga_com_tile_module_n_162, vga_com_tile_module_n_163 : std_logic;
  signal vga_com_tile_module_n_164, vga_com_tile_module_n_165, vga_com_tile_module_n_166, vga_com_tile_module_n_167, vga_com_tile_module_n_168 : std_logic;
  signal vga_com_tile_module_n_169, vga_com_tile_module_n_170, vga_com_tile_module_n_171, vga_com_tile_module_n_172, vga_com_tile_module_n_173 : std_logic;
  signal vga_com_tile_module_n_174, vga_com_tile_module_n_175, vga_com_tile_module_n_176, vga_com_tile_module_n_177, vga_com_tile_module_n_178 : std_logic;
  signal vga_com_tile_module_n_179, vga_com_tile_module_n_180, vga_com_tile_module_n_181, vga_com_tile_module_n_182, vga_com_tile_module_n_183 : std_logic;
  signal vga_com_tile_module_n_184, vga_com_tile_module_n_185, vga_com_tile_module_n_186, vga_com_tile_module_n_187, vga_com_tile_module_n_188 : std_logic;
  signal vga_com_tile_module_n_189, vga_com_tile_module_n_190, vga_com_tile_module_n_191, vga_com_tile_module_n_192, vga_com_tile_module_n_193 : std_logic;
  signal vga_com_tile_module_n_194, vga_com_tile_module_n_195, vga_com_tile_module_n_196, vga_com_tile_module_n_197, vga_com_tile_module_n_198 : std_logic;
  signal vga_com_tile_module_n_199, vga_com_tile_module_n_200, vga_com_tile_module_n_201, vga_com_tile_module_n_202, vga_com_tile_module_n_203 : std_logic;
  signal vga_com_tile_module_n_204, vga_com_tile_module_n_205, vga_com_tile_module_n_206, vga_com_tile_module_n_207, vga_com_tile_module_n_208 : std_logic;
  signal vga_com_tile_module_n_209, vga_com_tile_module_n_210, vga_com_tile_module_n_211, vga_com_tile_module_n_212, vga_com_tile_module_n_213 : std_logic;
  signal vga_com_tile_module_n_214, vga_com_tile_module_n_215, vga_com_tile_module_n_216, vga_com_tile_module_n_217, vga_com_tile_module_n_218 : std_logic;
  signal vga_com_tile_module_n_219, vga_com_tile_module_n_220, vga_com_tile_module_n_221, vga_com_tile_module_n_222, vga_com_tile_module_n_223 : std_logic;
  signal vga_com_tile_module_n_224, vga_com_tile_module_n_225, vga_com_tile_module_n_226, vga_com_tile_module_n_227, vga_com_tile_module_n_228 : std_logic;
  signal vga_com_tile_module_n_229, vga_com_tile_module_n_230, vga_com_tile_module_n_231, vga_com_tile_module_n_232, vga_com_tile_module_n_233 : std_logic;
  signal vga_com_tile_module_n_234, vga_com_tile_module_n_235, vga_com_tile_module_n_236, vga_com_tile_module_n_237, vga_com_tile_module_n_238 : std_logic;
  signal vga_com_tile_module_n_239, vga_com_tile_module_n_240, vga_com_tile_module_n_241, vga_com_tile_module_n_242, vga_com_tile_module_n_243 : std_logic;
  signal vga_com_tile_module_n_244, vga_com_tile_module_n_245, vga_com_tile_module_n_246, vga_com_tile_module_n_247, vga_com_tile_module_n_248 : std_logic;
  signal vga_com_tile_module_n_249, vga_com_tile_module_n_250, vga_com_tile_module_n_251, vga_com_tile_module_n_252, vga_com_tile_module_n_253 : std_logic;
  signal vga_com_tile_module_n_254, vga_com_tile_module_n_255, vga_com_tile_module_n_256, vga_com_tile_module_n_257, vga_com_tile_module_n_258 : std_logic;
  signal vga_com_tile_module_n_259, vga_com_tile_module_n_260, vga_com_tile_module_n_261, vga_com_tile_module_n_262, vga_com_tile_module_n_263 : std_logic;
  signal vga_com_tile_module_n_264, vga_com_tile_module_n_265, vga_com_tile_module_n_266, vga_com_tile_module_n_267, vga_com_tile_module_n_268 : std_logic;
  signal vga_com_tile_module_n_269, vga_com_tile_module_n_270, vga_com_tile_module_n_271, vga_com_tile_module_n_272, vga_com_tile_module_n_273 : std_logic;
  signal vga_com_tile_module_n_274, vga_com_tile_module_n_275, vga_com_tile_module_n_276, vga_com_tile_module_n_277, vga_com_tile_module_n_278 : std_logic;
  signal vga_com_tile_module_n_279, vga_com_tile_module_n_280, vga_com_tile_module_n_281, vga_com_tile_module_n_282, vga_com_tile_module_n_283 : std_logic;
  signal vga_com_tile_module_n_284, vga_com_tile_module_n_285, vga_com_tile_module_n_286, vga_com_tile_module_n_287, vga_com_tile_module_n_288 : std_logic;
  signal vga_com_tile_module_n_289, vga_com_tile_module_n_290, vga_com_tile_module_n_291, vga_com_tile_module_n_292, vga_com_tile_module_n_293 : std_logic;
  signal vga_com_tile_module_n_294, vga_com_tile_module_n_295, vga_com_tile_module_n_296, vga_com_tile_module_n_297, vga_com_tile_module_n_298 : std_logic;
  signal vga_com_tile_module_n_299, vga_com_tile_module_n_300, vga_com_tile_module_n_301, vga_com_tile_module_n_302, vga_com_tile_module_n_303 : std_logic;
  signal vga_com_tile_module_n_304, vga_com_tile_module_n_305, vga_com_tile_module_n_306, vga_com_tile_module_n_307, vga_com_tile_module_n_308 : std_logic;
  signal vga_com_tile_module_n_309, vga_com_tile_module_n_310, vga_com_tile_module_n_311, vga_com_tile_module_n_312, vga_com_tile_module_n_313 : std_logic;
  signal vga_com_tile_module_n_314, vga_com_tile_module_n_315, vga_com_tile_module_n_316, vga_com_tile_module_n_317, vga_com_tile_module_n_318 : std_logic;
  signal vga_com_tile_module_n_319, vga_com_tile_module_n_320, vga_com_tile_module_n_321, vga_com_tile_module_n_322, vga_com_tile_module_n_323 : std_logic;
  signal vga_com_tile_module_n_324, vga_com_tile_module_n_325, vga_com_tile_module_n_326, vga_com_tile_module_n_327, vga_com_tile_module_n_328 : std_logic;
  signal vga_com_tile_module_n_329, vga_com_tile_module_n_330, vga_com_tile_module_n_331, vga_com_tile_module_n_332, vga_com_tile_module_n_333 : std_logic;
  signal vga_com_tile_module_n_334, vga_com_tile_module_n_335, vga_com_tile_module_n_336, vga_com_tile_module_n_337, vga_com_tile_module_n_338 : std_logic;
  signal vga_com_tile_module_n_339, vga_com_tile_module_n_340, vga_com_tile_module_n_341, vga_com_tile_module_n_342, vga_com_tile_module_n_343 : std_logic;
  signal vga_com_tile_module_n_344, vga_com_tile_module_n_345, vga_com_tile_module_n_346, vga_com_tile_module_n_347, vga_com_tile_module_n_348 : std_logic;
  signal vga_com_tile_module_n_349, vga_com_tile_module_n_350, vga_com_tile_module_n_351, vga_com_tile_module_n_352, vga_com_tile_module_n_353 : std_logic;
  signal vga_com_tile_module_n_354, vga_com_tile_module_n_355, vga_com_tile_module_n_356, vga_com_tile_module_n_357, vga_com_tile_module_n_358 : std_logic;
  signal vga_com_tile_module_n_359, vga_com_tile_module_n_360, vga_com_tile_module_n_361, vga_com_tile_module_n_362, vga_com_tile_module_n_363 : std_logic;
  signal vga_com_tile_module_n_364, vga_com_tile_module_n_365, vga_com_tile_module_n_366, vga_com_tile_module_n_367, vga_com_tile_module_n_368 : std_logic;
  signal vga_com_tile_module_n_369, vga_com_tile_module_n_370, vga_com_tile_module_n_371, vga_com_tile_module_n_372, vga_com_tile_module_n_373 : std_logic;
  signal vga_com_tile_module_n_374, vga_com_tile_module_n_375, vga_com_tile_module_n_376, vga_com_tile_module_n_377, vga_com_tile_module_n_378 : std_logic;
  signal vga_com_tile_module_n_379, vga_com_tile_module_n_380, vga_com_tile_module_n_381, vga_com_tile_module_n_382, vga_com_tile_module_n_383 : std_logic;
  signal vga_com_tile_module_n_384, vga_com_tile_module_n_385, vga_com_tile_module_n_386, vga_com_tile_module_n_387, vga_com_tile_module_n_388 : std_logic;
  signal vga_com_tile_module_n_389, vga_com_tile_module_n_390, vga_com_tile_module_n_391, vga_com_tile_module_n_392, vga_com_tile_module_n_393 : std_logic;
  signal vga_com_tile_module_n_394, vga_com_tile_module_n_395, vga_com_tile_module_n_396, vga_com_tile_module_n_397, vga_com_tile_module_n_398 : std_logic;
  signal vga_com_tile_module_n_399, vga_com_tile_module_n_400, vga_com_tile_module_n_401, vga_com_tile_module_n_402, vga_com_tile_module_n_403 : std_logic;
  signal vga_com_tile_module_n_404, vga_com_tile_module_n_405, vga_com_tile_module_n_406, vga_com_tile_module_n_407, vga_com_tile_module_n_408 : std_logic;
  signal vga_com_tile_module_n_409, vga_com_tile_module_n_410, vga_com_tile_module_n_411, vga_com_tile_module_n_412, vga_com_tile_module_n_413 : std_logic;
  signal vga_com_tile_module_n_414, vga_com_tile_module_n_415, vga_com_tile_module_n_416, vga_com_tile_module_n_417, vga_com_tile_module_n_418 : std_logic;
  signal vga_com_tile_module_n_419, vga_com_tile_module_n_420, vga_com_tile_module_n_421, vga_com_tile_module_n_422, vga_com_tile_module_n_423 : std_logic;
  signal vga_com_tile_module_n_424, vga_com_tile_module_n_425, vga_com_tile_module_n_426, vga_com_tile_module_n_427, vga_com_tile_module_n_428 : std_logic;
  signal vga_com_tile_module_n_429, vga_com_tile_module_n_430, vga_com_tile_module_n_431, vga_com_tile_module_n_432, vga_com_tile_module_n_433 : std_logic;
  signal vga_com_tile_module_n_434, vga_com_tile_module_n_435, vga_com_tile_module_n_436, vga_com_tile_module_n_437, vga_com_tile_module_n_438 : std_logic;
  signal vga_com_tile_module_n_439, vga_com_tile_module_n_440, vga_com_tile_module_n_441, vga_com_tile_module_n_442, vga_com_tile_module_n_443 : std_logic;
  signal vga_com_tile_module_n_444, vga_com_tile_module_n_445, vga_com_tile_module_n_446, vga_com_tile_module_n_447, vga_com_tile_module_n_448 : std_logic;
  signal vga_com_tile_module_n_449, vga_com_tile_module_n_450, vga_com_tile_module_n_451, vga_com_tile_module_n_452, vga_com_tile_module_n_453 : std_logic;
  signal vga_com_tile_module_n_454, vga_com_tile_module_n_455, vga_com_tile_module_n_456, vga_com_tile_module_n_457, vga_com_tile_module_n_458 : std_logic;
  signal vga_com_tile_module_n_459, vga_com_tile_module_n_460, vga_com_tile_module_n_461, vga_com_tile_module_n_462, vga_com_tile_module_n_463 : std_logic;
  signal vga_com_tile_module_n_464, vga_com_tile_module_n_465, vga_com_tile_module_n_466, vga_com_tile_module_n_467, vga_com_tile_module_n_468 : std_logic;
  signal vga_com_tile_module_n_469, vga_com_tile_module_n_470, vga_com_tile_module_n_471, vga_com_tile_module_n_472, vga_com_tile_module_n_473 : std_logic;
  signal vga_com_tile_module_n_474, vga_com_tile_module_n_475, vga_com_tile_module_n_476, vga_com_tile_module_n_477, vga_com_tile_module_n_478 : std_logic;
  signal vga_com_tile_module_n_479, vga_com_tile_module_n_480, vga_com_tile_module_n_481, vga_com_tile_module_n_482, vga_com_tile_module_n_483 : std_logic;
  signal vga_com_tile_module_n_484, vga_com_tile_module_n_485, vga_com_tile_module_n_486, vga_com_tile_module_n_487, vga_com_tile_module_n_488 : std_logic;
  signal vga_com_tile_module_n_489, vga_com_tile_module_n_490, vga_com_tile_module_n_491, vga_com_tile_module_n_492, vga_com_tile_module_n_493 : std_logic;
  signal vga_com_tile_module_n_494, vga_com_tile_module_n_495, vga_com_tile_module_n_496, vga_com_tile_module_n_497, vga_com_tile_module_n_498 : std_logic;
  signal vga_com_tile_module_n_499, vga_com_tile_module_n_500, vga_com_tile_module_n_501, vga_com_tile_module_n_502, vga_com_tile_module_n_503 : std_logic;
  signal vga_com_tile_module_n_504, vga_com_tile_module_n_505, vga_com_tile_module_n_506, vga_com_tile_module_n_507, vga_com_tile_module_n_508 : std_logic;
  signal vga_com_tile_module_n_509, vga_com_tile_module_n_510, vga_com_tile_module_n_511, vga_com_tile_module_n_512, vga_com_tile_module_n_513 : std_logic;
  signal vga_com_tile_module_n_514, vga_com_tile_module_n_515, vga_com_tile_module_n_516, vga_com_tile_module_n_517, vga_com_tile_module_n_518 : std_logic;
  signal vga_com_tile_module_n_519, vga_com_tile_module_n_520, vga_com_tile_module_n_521, vga_com_tile_module_n_522, vga_com_tile_module_n_523 : std_logic;
  signal vga_com_tile_module_n_524, vga_com_tile_module_n_525, vga_com_tile_module_n_526, vga_com_tile_module_n_528, vga_com_tile_module_n_529 : std_logic;
  signal vga_com_tile_module_n_530, vga_com_tile_module_n_531, vga_com_tile_module_n_532, vga_com_tile_module_n_533, vga_com_tile_module_n_534 : std_logic;
  signal vga_com_tile_module_n_535, vga_com_tile_module_n_536, vga_com_tile_module_n_537, vga_com_tile_module_n_538, vga_com_tile_module_n_539 : std_logic;
  signal vga_com_tile_module_n_540, vga_com_tile_module_n_541, vga_com_tile_module_n_542, vga_com_tile_module_n_543, vga_com_tile_module_n_544 : std_logic;
  signal vga_com_tile_module_n_545, vga_com_tile_module_n_546, vga_com_tile_module_n_547, vga_com_tile_module_n_548, vga_com_tile_module_n_549 : std_logic;
  signal vga_com_tile_module_n_550, vga_com_tile_module_n_551, vga_com_tile_module_n_552, vga_com_tile_module_n_553, vga_com_tile_module_n_554 : std_logic;
  signal vga_com_tile_module_n_555, vga_com_tile_module_n_556, vga_com_tile_module_n_557, vga_com_tile_module_n_558, vga_com_tile_module_n_559 : std_logic;
  signal vga_com_tile_module_n_560, vga_com_tile_module_n_561, vga_com_tile_module_n_562, vga_com_tile_module_n_563, vga_com_tile_module_n_564 : std_logic;
  signal vga_com_tile_module_n_565, vga_com_tile_module_n_566, vga_com_tile_module_n_567, vga_com_tile_module_n_568, vga_com_tile_module_n_569 : std_logic;
  signal vga_com_tile_module_n_570, vga_com_tile_module_n_571, vga_com_tile_module_n_572, vga_com_tile_module_n_573, vga_com_tile_module_n_574 : std_logic;
  signal vga_com_tile_module_n_575, vga_com_tile_module_n_576, vga_com_tile_module_n_577, vga_com_tile_module_n_578, vga_com_tile_module_n_579 : std_logic;
  signal vga_com_tile_module_n_580, vga_com_tile_module_n_581, vga_com_tile_module_n_582, vga_com_tile_module_n_583, vga_com_tile_module_n_584 : std_logic;
  signal vga_com_tile_module_n_585, vga_com_tile_module_n_586, vga_com_tile_module_n_587, vga_com_tile_module_n_588, vga_com_tile_module_n_589 : std_logic;
  signal vga_com_tile_module_n_590, vga_com_tile_module_n_591, vga_com_tile_module_n_592, vga_com_tile_module_n_593, vga_com_tile_module_n_594 : std_logic;
  signal vga_com_tile_module_n_595, vga_com_tile_module_n_596, vga_com_tile_module_n_597, vga_com_tile_module_n_598, vga_com_tile_module_n_599 : std_logic;
  signal vga_com_tile_module_n_600, vga_com_tile_module_n_601, vga_com_tile_module_n_602, vga_com_tile_module_n_603, vga_com_tile_module_n_604 : std_logic;
  signal vga_com_tile_module_n_605, vga_com_tile_module_n_606, vga_com_tile_module_n_607, vga_com_tile_module_n_608, vga_com_tile_module_n_609 : std_logic;
  signal vga_com_tile_module_n_610, vga_com_tile_module_n_611, vga_com_tile_module_n_612, vga_com_tile_module_n_613, vga_com_tile_module_n_614 : std_logic;
  signal vga_com_tile_module_n_615, vga_com_tile_module_n_616, vga_com_tile_module_n_617, vga_com_tile_module_n_618, vga_com_tile_module_n_619 : std_logic;
  signal vga_com_tile_module_n_620, vga_com_tile_module_n_621, vga_com_tile_module_n_622, vga_com_tile_module_n_623, vga_com_tile_module_n_624 : std_logic;
  signal vga_com_tile_module_n_625, vga_com_tile_module_n_626, vga_com_tile_module_n_627, vga_com_tile_module_n_628, vga_com_tile_module_n_629 : std_logic;
  signal vga_com_tile_module_n_630, vga_com_tile_module_n_631, vga_com_tile_module_n_632, vga_com_tile_module_n_633, vga_com_tile_module_n_634 : std_logic;
  signal vga_com_tile_module_n_635, vga_com_tile_module_n_636, vga_com_tile_module_n_637, vga_com_tile_module_n_638, vga_com_tile_module_n_639 : std_logic;
  signal vga_com_tile_module_n_640, vga_com_tile_module_n_641, vga_com_tile_module_n_642, vga_com_tile_module_n_643, vga_com_tile_module_n_644 : std_logic;
  signal vga_com_tile_module_n_645, vga_com_tile_module_n_646, vga_com_tile_module_n_647, vga_com_tile_module_n_648, vga_com_tile_module_n_649 : std_logic;
  signal vga_com_tile_module_n_650, vga_com_tile_module_n_651, vga_com_tile_module_n_652, vga_com_tile_module_n_653, vga_com_tile_module_n_654 : std_logic;
  signal vga_com_tile_module_n_655, vga_com_tile_module_n_656, vga_com_tile_module_n_657, vga_com_tile_module_n_658, vga_com_tile_module_n_659 : std_logic;
  signal vga_com_tile_module_n_660, vga_com_tile_module_n_661, vga_com_tile_module_n_662, vga_com_tile_module_n_663, vga_com_tile_module_n_664 : std_logic;
  signal vga_com_tile_module_n_665, vga_com_tile_module_n_666, vga_com_tile_module_n_667, vga_com_tile_module_n_668, vga_com_tile_module_n_669 : std_logic;
  signal vga_com_tile_module_n_670, vga_com_tile_module_n_671, vga_com_tile_module_n_672, vga_com_tile_module_n_673, vga_com_tile_module_n_674 : std_logic;
  signal vga_com_tile_module_n_675, vga_com_tile_module_n_676, vga_com_tile_module_n_677, vga_com_tile_module_n_678, vga_com_tile_module_n_679 : std_logic;
  signal vga_com_tile_module_n_680, vga_com_tile_module_n_681, vga_com_tile_module_n_682, vga_com_tile_module_n_683, vga_com_tile_module_n_684 : std_logic;
  signal vga_com_tile_module_n_685, vga_com_tile_module_n_686, vga_com_tile_module_n_687, vga_com_tile_module_n_688, vga_com_tile_module_n_689 : std_logic;
  signal vga_com_tile_module_n_690, vga_com_tile_module_n_691, vga_com_tile_module_n_692, vga_com_tile_module_n_693, vga_com_tile_module_n_694 : std_logic;
  signal vga_com_tile_module_n_695, vga_com_tile_module_n_696, vga_com_tile_module_n_697, vga_com_tile_module_n_698, vga_com_tile_module_n_699 : std_logic;
  signal vga_com_tile_module_n_700, vga_com_tile_module_n_701, vga_com_tile_module_n_702, vga_com_tile_module_n_703, vga_com_tile_module_n_704 : std_logic;
  signal vga_com_tile_module_n_705, vga_com_tile_module_n_706, vga_com_tile_module_n_707, vga_com_tile_module_n_708, vga_com_tile_module_n_709 : std_logic;
  signal vga_com_tile_module_n_710, vga_com_tile_module_n_711, vga_com_tile_module_n_712, vga_com_tile_module_n_713, vga_com_tile_module_n_714 : std_logic;
  signal vga_com_tile_module_n_715, vga_com_tile_module_n_716, vga_com_tile_module_n_717, vga_com_tile_module_n_718, vga_com_tile_module_n_719 : std_logic;
  signal vga_com_tile_module_n_720, vga_com_tile_module_n_721, vga_com_tile_module_n_722, vga_com_tile_module_n_723, vga_com_tile_module_n_724 : std_logic;
  signal vga_com_tile_module_n_725, vga_com_tile_module_n_726, vga_com_tile_module_n_727, vga_com_tile_module_n_728, vga_com_tile_module_n_729 : std_logic;
  signal vga_com_tile_module_n_730, vga_com_tile_module_n_731, vga_com_tile_module_n_732, vga_com_tile_module_n_733, vga_com_tile_module_n_734 : std_logic;
  signal vga_com_tile_module_n_735, vga_com_tile_module_n_736, vga_com_tile_module_n_737, vga_com_tile_module_n_738, vga_com_tile_module_n_739 : std_logic;
  signal vga_com_tile_module_n_740, vga_com_tile_module_n_741, vga_com_tile_module_n_742, vga_com_tile_module_n_743, vga_com_tile_module_n_744 : std_logic;
  signal vga_com_tile_module_n_745, vga_com_tile_module_n_746, vga_com_tile_module_n_747, vga_com_tile_module_n_748, vga_com_tile_module_n_749 : std_logic;
  signal vga_com_tile_module_n_750, vga_com_tile_module_n_751, vga_com_tile_module_n_752, vga_com_tile_module_n_753, vga_com_tile_module_n_754 : std_logic;
  signal vga_com_tile_module_n_755, vga_com_tile_module_n_756, vga_com_tile_module_n_757, vga_com_tile_module_n_758, vga_com_tile_module_n_759 : std_logic;
  signal vga_com_tile_module_n_760, vga_com_tile_module_n_761, vga_com_tile_module_n_762, vga_com_tile_module_n_763, vga_com_tile_module_n_764 : std_logic;
  signal vga_com_tile_module_n_765, vga_com_tile_module_n_766, vga_com_tile_module_n_767, vga_com_tile_module_n_768, vga_com_tile_module_n_769 : std_logic;
  signal vga_com_tile_module_n_770, vga_com_tile_module_n_771, vga_com_tile_module_n_772, vga_com_tile_module_n_773, vga_com_tile_module_n_774 : std_logic;
  signal vga_com_tile_module_n_775, vga_com_tile_module_n_776, vga_com_tile_module_n_777, vga_com_tile_module_n_778, vga_com_tile_module_n_779 : std_logic;
  signal vga_com_tile_module_n_780, vga_com_tile_module_n_781, vga_com_tile_module_n_782, vga_com_tile_module_n_783, vga_com_tile_module_n_784 : std_logic;
  signal vga_com_tile_module_n_785, vga_com_tile_module_n_786, vga_com_tile_module_n_787, vga_com_tile_module_n_788, vga_com_tile_module_n_789 : std_logic;
  signal vga_com_tile_module_n_790, vga_com_tile_module_n_791, vga_com_tile_module_n_792, vga_com_tile_module_n_793, vga_com_tile_module_n_794 : std_logic;
  signal vga_com_tile_module_n_795, vga_com_tile_module_n_796, vga_com_tile_module_n_797, vga_com_tile_module_n_798, vga_com_tile_module_n_799 : std_logic;
  signal vga_com_tile_module_n_800, vga_com_tile_module_n_801, vga_com_tile_module_n_802, vga_com_tile_module_n_803, vga_com_tile_module_n_804 : std_logic;
  signal vga_com_tile_module_n_805, vga_com_tile_module_n_806, vga_com_tile_module_n_807, vga_com_tile_module_n_808, vga_com_tile_module_n_809 : std_logic;
  signal vga_com_tile_module_n_810, vga_com_tile_module_n_811, vga_com_tile_module_n_812, vga_com_tile_module_n_813, vga_com_tile_module_n_814 : std_logic;
  signal vga_com_tile_module_n_815, vga_com_tile_module_n_816, vga_com_tile_module_n_817, vga_com_tile_module_n_818, vga_com_tile_module_n_819 : std_logic;
  signal vga_com_tile_module_n_820, vga_com_tile_module_n_821, vga_com_tile_module_n_822, vga_com_tile_module_n_823, vga_com_tile_module_n_824 : std_logic;
  signal vga_com_tile_module_n_825, vga_com_tile_module_n_826, vga_com_tile_module_n_827, vga_com_tile_module_n_828, vga_com_tile_module_n_829 : std_logic;
  signal vga_com_tile_module_n_830, vga_com_tile_module_n_831, vga_com_tile_module_n_832, vga_com_tile_module_n_833, vga_com_tile_module_n_834 : std_logic;
  signal vga_com_tile_module_n_835, vga_com_tile_module_n_836, vga_com_tile_module_n_837, vga_com_tile_module_n_838, vga_com_tile_module_n_839 : std_logic;
  signal vga_com_tile_module_n_840, vga_com_tile_module_n_841, vga_com_tile_module_n_842, vga_com_tile_module_n_843, vga_com_tile_module_n_844 : std_logic;
  signal vga_com_tile_module_n_845, vga_com_tile_module_n_846, vga_com_tile_module_n_847, vga_com_tile_module_n_848, vga_com_tile_module_n_849 : std_logic;
  signal vga_com_tile_module_n_850, vga_com_tile_module_n_851, vga_com_tile_module_n_852, vga_com_tile_module_n_853, vga_com_tile_module_n_854 : std_logic;
  signal vga_com_tile_module_n_855, vga_com_tile_module_n_856, vga_com_tile_module_n_857, vga_com_tile_module_n_858, vga_com_tile_module_n_859 : std_logic;
  signal vga_com_tile_module_n_860, vga_com_tile_module_n_861, vga_com_tile_module_n_862, vga_com_tile_module_n_863, vga_com_tile_module_n_864 : std_logic;
  signal vga_com_tile_module_n_865, vga_com_tile_module_n_866, vga_com_tile_module_n_867, vga_com_tile_module_n_868, vga_com_tile_module_n_869 : std_logic;
  signal vga_com_tile_module_n_870, vga_com_tile_module_n_871, vga_com_tile_module_n_872, vga_com_tile_module_n_873, vga_com_tile_module_n_874 : std_logic;
  signal vga_com_tile_module_n_875, vga_com_tile_module_n_876, vga_com_tile_module_n_877, vga_com_tile_module_n_878, vga_com_tile_module_n_879 : std_logic;
  signal vga_com_tile_module_n_880, vga_com_tile_module_n_881, vga_com_tile_module_n_882, vga_com_tile_module_n_883, vga_com_tile_module_n_884 : std_logic;
  signal vga_com_tile_module_n_885, vga_com_tile_module_n_886, vga_com_tile_module_n_887, vga_com_tile_module_n_888, vga_com_tile_module_n_889 : std_logic;
  signal vga_com_tile_module_n_890, vga_com_tile_module_n_891, vga_com_tile_module_n_892, vga_com_tile_module_n_893, vga_com_tile_module_n_894 : std_logic;
  signal vga_com_tile_module_n_895, vga_com_tile_module_n_896, vga_com_tile_module_n_897, vga_com_tile_module_n_898, vga_com_tile_module_n_899 : std_logic;
  signal vga_com_tile_module_n_900, vga_com_tile_module_n_901, vga_com_tile_module_n_902, vga_com_tile_module_n_903, vga_com_tile_module_n_904 : std_logic;
  signal vga_com_tile_module_n_905, vga_com_tile_module_n_906, vga_com_tile_module_n_907, vga_com_tile_module_n_908, vga_com_tile_module_n_909 : std_logic;
  signal vga_com_tile_module_n_910, vga_com_tile_module_n_911, vga_com_tile_module_n_912, vga_com_tile_module_n_913, vga_com_tile_module_n_914 : std_logic;
  signal vga_com_tile_module_n_915, vga_com_tile_module_n_916, vga_com_tile_module_n_917, vga_com_tile_module_n_918, vga_com_tile_module_n_919 : std_logic;
  signal vga_com_tile_module_n_920, vga_com_tile_module_n_921, vga_com_tile_module_n_922, vga_com_tile_module_n_923, vga_com_tile_module_n_924 : std_logic;
  signal vga_com_tile_module_n_925, vga_com_tile_module_n_926, vga_com_tile_module_n_927, vga_com_tile_module_n_928, vga_com_tile_module_n_929 : std_logic;
  signal vga_com_tile_module_n_930, vga_com_tile_module_n_931, vga_com_tile_module_n_932, vga_com_tile_module_n_933, vga_com_tile_module_n_934 : std_logic;
  signal vga_com_tile_module_n_935, vga_com_tile_module_n_936, vga_com_tile_module_n_937, vga_com_tile_module_n_938, vga_com_tile_module_n_939 : std_logic;
  signal vga_com_tile_module_n_940, vga_com_tile_module_n_941, vga_com_tile_module_n_942, vga_com_tile_module_n_943, vga_com_tile_module_n_944 : std_logic;
  signal vga_com_tile_module_n_945, vga_com_tile_module_n_946, vga_com_tile_module_n_947, vga_com_tile_module_n_948, vga_com_tile_module_n_949 : std_logic;
  signal vga_com_tile_module_n_950, vga_com_tile_module_n_951, vga_com_tile_module_n_952, vga_com_tile_module_n_953, vga_com_tile_module_n_954 : std_logic;
  signal vga_com_tile_module_n_955, vga_com_tile_module_n_956, vga_com_tile_module_n_957, vga_com_tile_module_n_958, vga_com_tile_module_n_959 : std_logic;
  signal vga_com_tile_module_n_960, vga_com_tile_module_n_961, vga_com_tile_module_n_962, vga_com_tile_module_n_963, vga_com_tile_module_n_964 : std_logic;
  signal vga_com_tile_module_n_965, vga_com_tile_module_n_966, vga_com_tile_module_n_967, vga_com_tile_module_n_968, vga_com_tile_module_n_969 : std_logic;
  signal vga_com_tile_module_n_970, vga_com_tile_module_n_971, vga_com_tile_module_n_972, vga_com_tile_module_n_973, vga_com_tile_module_n_974 : std_logic;
  signal vga_com_tile_module_n_975, vga_com_tile_module_n_976, vga_com_tile_module_n_977, vga_com_tile_module_n_978, vga_com_tile_module_n_979 : std_logic;
  signal vga_com_tile_module_n_980, vga_com_tile_module_n_981, vga_com_tile_module_n_982, vga_com_tile_module_n_983, vga_com_tile_module_n_984 : std_logic;
  signal vga_com_tile_module_n_985, vga_com_tile_module_n_986, vga_com_tile_module_n_987, vga_com_tile_module_n_988, vga_com_tile_module_n_989 : std_logic;
  signal vga_com_tile_module_n_990, vga_com_tile_module_n_991, vga_com_tile_module_n_992, vga_com_tile_module_n_993, vga_com_tile_module_n_994 : std_logic;
  signal vga_com_tile_module_n_995, vga_com_tile_module_n_996, vga_com_tile_module_n_997, vga_com_tile_module_n_998, vga_com_tile_module_n_999 : std_logic;
  signal vga_com_tile_module_n_1000, vga_com_tile_module_n_1001, vga_com_tile_module_n_1002, vga_com_tile_module_n_1003, vga_com_tile_module_n_1004 : std_logic;
  signal vga_com_tile_module_n_1005, vga_com_tile_module_n_1006, vga_com_tile_module_n_1007, vga_com_tile_module_n_1008, vga_com_tile_module_n_1009 : std_logic;
  signal vga_com_tile_module_n_1010, vga_com_tile_module_n_1011, vga_com_tile_module_n_1012, vga_com_tile_module_n_1013, vga_com_tile_module_n_1014 : std_logic;
  signal vga_com_tile_module_n_1015, vga_com_tile_module_n_1016, vga_com_tile_module_n_1017, vga_com_tile_module_n_1018, vga_com_tile_module_n_1019 : std_logic;
  signal vga_com_tile_module_n_1020, vga_com_tile_module_n_1021, vga_com_tile_module_n_1022, vga_com_tile_module_n_1023, vga_com_tile_module_n_1024 : std_logic;
  signal vga_com_tile_module_n_1025, vga_com_tile_module_n_1026, vga_com_tile_module_n_1027, vga_com_tile_module_n_1028, vga_com_tile_module_n_1029 : std_logic;
  signal vga_com_tile_module_n_1030, vga_com_tile_module_n_1031, vga_com_tile_module_n_1033, vga_com_tile_module_n_1034, vga_com_tile_module_n_1038 : std_logic;
  signal vga_com_tile_module_n_1039, vga_com_tile_module_n_1040, vga_com_tile_module_n_1041, vga_com_tile_module_n_1060, vga_done : std_logic;

begin

  FE_PHC510_map_data_9 : BUFFD2BWP7T port map(I => FE_PHN425_map_data_9, Z => FE_PHN510_map_data_9);
  FE_PHC509_map_data_56 : BUFFD2BWP7T port map(I => FE_PHN509_map_data_56, Z => map_data(56));
  FE_PHC508_stable_map_com_n_86 : BUFFD2BWP7T port map(I => stable_map_com_n_86, Z => FE_PHN508_stable_map_com_n_86);
  FE_PHC507_map_data_24 : BUFFD1P5BWP7T port map(I => map_data(24), Z => FE_PHN507_map_data_24);
  FE_PHC506_map_data_30 : DEL01BWP7T port map(I => FE_PHN506_map_data_30, Z => map_data(30));
  FE_PHC505_map_data_42 : BUFFD1P5BWP7T port map(I => map_data(42), Z => FE_PHN505_map_data_42);
  FE_PHC504_map_data_26 : BUFFD1P5BWP7T port map(I => FE_PHN501_map_data_26, Z => FE_PHN504_map_data_26);
  FE_PHC503_map_data_40 : BUFFD1P5BWP7T port map(I => map_data(40), Z => FE_PHN503_map_data_40);
  FE_PHC502_fsm_com_n_489 : DEL01BWP7T port map(I => FE_PHN487_fsm_com_n_489, Z => FE_PHN502_fsm_com_n_489);
  FE_PHC501_map_data_26 : CKBD2BWP7T port map(I => map_data(26), Z => FE_PHN501_map_data_26);
  FE_PHC500_map_data_16 : BUFFD2BWP7T port map(I => FE_PHN481_map_data_16, Z => FE_PHN500_map_data_16);
  FE_PHC499_map_data_32 : BUFFD2BWP7T port map(I => FE_PHN474_map_data_32, Z => FE_PHN499_map_data_32);
  FE_PHC498_level_d_1 : DEL01BWP7T port map(I => FE_PHN454_level_d_1, Z => FE_PHN498_level_d_1);
  FE_PHC497_map_data_22 : BUFFD2BWP7T port map(I => map_data(22), Z => FE_PHN497_map_data_22);
  FE_PHC496_map_data_15 : BUFFD2BWP7T port map(I => FE_PHN475_map_data_15, Z => FE_PHN496_map_data_15);
  FE_PHC495_map_data_45 : BUFFD2BWP7T port map(I => map_data(45), Z => FE_PHN495_map_data_45);
  FE_PHC494_spi_com_n_74 : DEL01BWP7T port map(I => FE_PHN479_spi_com_n_74, Z => FE_PHN494_spi_com_n_74);
  FE_PHC493_map_data_25 : BUFFD0BWP7T port map(I => FE_PHN435_map_data_25, Z => FE_PHN493_map_data_25);
  FE_PHC492_stable_map_com_n_79 : DEL01BWP7T port map(I => FE_PHN488_stable_map_com_n_79, Z => FE_PHN492_stable_map_com_n_79);
  FE_PHC491_map_data_29 : CKBD2BWP7T port map(I => FE_PHN437_map_data_29, Z => FE_PHN491_map_data_29);
  FE_PHC490_map_data_31 : BUFFD0BWP7T port map(I => map_data(31), Z => FE_PHN490_map_data_31);
  FE_PHC489_level_d_1 : CKBD0BWP7T port map(I => level_d(1), Z => FE_PHN489_level_d_1);
  FE_PHC488_stable_map_com_n_79 : CKBD0BWP7T port map(I => FE_PHN433_stable_map_com_n_79, Z => FE_PHN488_stable_map_com_n_79);
  FE_PHC487_fsm_com_n_489 : CKBD0BWP7T port map(I => FE_PHN459_fsm_com_n_489, Z => FE_PHN487_fsm_com_n_489);
  FE_PHC486_map_data_28 : CKBD0BWP7T port map(I => FE_PHN449_map_data_28, Z => FE_PHN486_map_data_28);
  FE_PHC485_map_data_55 : CKBD0BWP7T port map(I => FE_PHN428_map_data_55, Z => FE_PHN485_map_data_55);
  FE_PHC484_map_data_47 : CKBD0BWP7T port map(I => FE_PHN444_map_data_47, Z => FE_PHN484_map_data_47);
  FE_PHC483_map_data_59 : CKBD0BWP7T port map(I => FE_PHN451_map_data_59, Z => FE_PHN483_map_data_59);
  FE_PHC482_map_data_30 : CKBD0BWP7T port map(I => FE_PHN447_map_data_30, Z => FE_PHN482_map_data_30);
  FE_PHC481_map_data_16 : CKBD0BWP7T port map(I => FE_PHN450_map_data_16, Z => FE_PHN481_map_data_16);
  FE_PHC480_map_data_56 : CKBD0BWP7T port map(I => FE_PHN429_map_data_56, Z => FE_PHN480_map_data_56);
  FE_PHC479_spi_com_n_74 : CKBD0BWP7T port map(I => FE_PHN420_spi_com_n_74, Z => FE_PHN479_spi_com_n_74);
  FE_PHC478_map_data_50 : CKBD0BWP7T port map(I => FE_PHN452_map_data_50, Z => FE_PHN478_map_data_50);
  FE_PHC477_level_d_4 : DEL01BWP7T port map(I => FE_PHN413_level_d_4, Z => FE_PHN477_level_d_4);
  FE_PHC476_map_data_21 : CKBD0BWP7T port map(I => FE_PHN424_map_data_21, Z => FE_PHN476_map_data_21);
  FE_PHC475_map_data_15 : CKBD0BWP7T port map(I => FE_PHN431_map_data_15, Z => FE_PHN475_map_data_15);
  FE_PHC474_map_data_32 : CKBD0BWP7T port map(I => FE_PHN446_map_data_32, Z => FE_PHN474_map_data_32);
  FE_PHC473_map_data_39 : CKBD0BWP7T port map(I => FE_PHN434_map_data_39, Z => FE_PHN473_map_data_39);
  FE_PHC472_map_data_60 : CKBD0BWP7T port map(I => FE_PHN448_map_data_60, Z => FE_PHN472_map_data_60);
  FE_PHC471_stable_map_com_n_84 : DEL01BWP7T port map(I => FE_PHN412_stable_map_com_n_84, Z => FE_PHN471_stable_map_com_n_84);
  FE_PHC470_map_data_41 : CKBD0BWP7T port map(I => FE_PHN422_map_data_41, Z => FE_PHN470_map_data_41);
  FE_PHC469_map_data_45 : CKBD0BWP7T port map(I => FE_PHN436_map_data_45, Z => FE_PHN469_map_data_45);
  FE_PHC468_map_data_43 : CKBD0BWP7T port map(I => FE_PHN443_map_data_43, Z => FE_PHN468_map_data_43);
  FE_PHC467_map_data_22 : CKBD0BWP7T port map(I => FE_PHN442_map_data_22, Z => FE_PHN467_map_data_22);
  FE_PHC466_map_data_40 : CKBD0BWP7T port map(I => FE_PHN445_map_data_40, Z => FE_PHN466_map_data_40);
  FE_PHC465_map_data_4 : DEL01BWP7T port map(I => map_data(4), Z => FE_PHN465_map_data_4);
  FE_PHC464_map_data_24 : CKBD0BWP7T port map(I => FE_PHN432_map_data_24, Z => FE_PHN464_map_data_24);
  FE_PHC463_map_data_42 : DEL02BWP7T port map(I => FE_PHN505_map_data_42, Z => FE_PHN463_map_data_42);
  FE_PHC462_spi_com_MISO_shift_42 : DEL01BWP7T port map(I => FE_PHN462_spi_com_MISO_shift_42, Z => FE_PHN366_spi_com_MISO_shift_42);
  FE_PHC461_map_data_8 : CKBD0BWP7T port map(I => FE_PHN417_map_data_8, Z => FE_PHN461_map_data_8);
  FE_PHC460_stable_map_com_n_102 : CKBD0BWP7T port map(I => FE_PHN460_stable_map_com_n_102, Z => FE_PHN430_stable_map_com_n_102);
  FE_PHC459_fsm_com_n_489 : CKBD0BWP7T port map(I => fsm_com_n_489, Z => FE_PHN459_fsm_com_n_489);
  FE_PHC458_energy_d_7 : DEL01BWP7T port map(I => FE_PHN458_energy_d_7, Z => energy_d(7));
  FE_PHC457_map_data_64 : DEL02BWP7T port map(I => FE_PHN457_map_data_64, Z => map_data(64));
  FE_PHC456_fsm_com_energy_8 : DEL01BWP7T port map(I => fsm_com_energy(8), Z => FE_PHN456_fsm_com_energy_8);
  FE_PHC455_spi_com_MISO_shift_42 : DEL015BWP7T port map(I => spi_com_MISO_shift(42), Z => FE_PHN455_spi_com_MISO_shift_42);
  FE_PHC454_level_d_1 : DEL02BWP7T port map(I => FE_PHN489_level_d_1, Z => FE_PHN454_level_d_1);
  FE_PHC453_spi_com_MISO_shift_34 : BUFFD1P5BWP7T port map(I => FE_PHN453_spi_com_MISO_shift_34, Z => FE_PHN369_spi_com_MISO_shift_34);
  FE_PHC452_map_data_50 : CKBD0BWP7T port map(I => map_data(50), Z => FE_PHN452_map_data_50);
  FE_PHC451_map_data_59 : CKBD0BWP7T port map(I => map_data(59), Z => FE_PHN451_map_data_59);
  FE_PHC450_map_data_16 : CKBD0BWP7T port map(I => map_data(16), Z => FE_PHN450_map_data_16);
  FE_PHC449_map_data_28 : CKBD0BWP7T port map(I => map_data(28), Z => FE_PHN449_map_data_28);
  FE_PHC448_map_data_60 : CKBD0BWP7T port map(I => map_data(60), Z => FE_PHN448_map_data_60);
  FE_PHC447_map_data_30 : CKBD0BWP7T port map(I => map_data(30), Z => FE_PHN447_map_data_30);
  FE_PHC446_map_data_32 : CKBD0BWP7T port map(I => map_data(32), Z => FE_PHN446_map_data_32);
  FE_PHC445_map_data_40 : CKBD0BWP7T port map(I => FE_PHN503_map_data_40, Z => FE_PHN445_map_data_40);
  FE_PHC444_map_data_47 : CKBD0BWP7T port map(I => map_data(47), Z => FE_PHN444_map_data_47);
  FE_PHC443_map_data_43 : CKBD0BWP7T port map(I => map_data(43), Z => FE_PHN443_map_data_43);
  FE_PHC442_map_data_22 : CKBD0BWP7T port map(I => FE_PHN497_map_data_22, Z => FE_PHN442_map_data_22);
  FE_PHC441_spi_com_MISO_shift_14 : DEL01BWP7T port map(I => FE_PHN190_spi_com_MISO_shift_14, Z => FE_PHN441_spi_com_MISO_shift_14);
  FE_PHC440_map_data_31 : CKBD2BWP7T port map(I => FE_PHN490_map_data_31, Z => FE_PHN440_map_data_31);
  FE_PHC439_map_data_11 : CKBD2BWP7T port map(I => map_data(11), Z => FE_PHN439_map_data_11);
  FE_PHC438_map_data_3 : CKBD2BWP7T port map(I => map_data(3), Z => FE_PHN438_map_data_3);
  FE_PHC437_map_data_29 : CKBD0BWP7T port map(I => map_data(29), Z => FE_PHN437_map_data_29);
  FE_PHC436_map_data_45 : BUFFD0BWP7T port map(I => FE_PHN495_map_data_45, Z => FE_PHN436_map_data_45);
  FE_PHC435_map_data_25 : BUFFD0BWP7T port map(I => map_data(25), Z => FE_PHN435_map_data_25);
  FE_PHC434_map_data_39 : CKBD0BWP7T port map(I => map_data(39), Z => FE_PHN434_map_data_39);
  FE_PHC433_stable_map_com_n_79 : CKBD0BWP7T port map(I => stable_map_com_n_79, Z => FE_PHN433_stable_map_com_n_79);
  FE_PHC432_map_data_24 : CKBD0BWP7T port map(I => FE_PHN507_map_data_24, Z => FE_PHN432_map_data_24);
  FE_PHC431_map_data_15 : CKBD0BWP7T port map(I => map_data(15), Z => FE_PHN431_map_data_15);
  FE_PHC430_stable_map_com_n_102 : CKBD0BWP7T port map(I => FE_PHN430_stable_map_com_n_102, Z => stable_map_com_n_102);
  FE_PHC429_map_data_56 : CKBD0BWP7T port map(I => map_data(56), Z => FE_PHN429_map_data_56);
  FE_PHC428_map_data_55 : CKBD0BWP7T port map(I => map_data(55), Z => FE_PHN428_map_data_55);
  FE_PHC427_stable_map_com_n_58 : CKBD0BWP7T port map(I => stable_map_com_n_58, Z => FE_PHN427_stable_map_com_n_58);
  FE_PHC426_map_data_42 : CKBD0BWP7T port map(I => FE_PHN463_map_data_42, Z => FE_PHN426_map_data_42);
  FE_PHC425_map_data_9 : CKBD0BWP7T port map(I => map_data(9), Z => FE_PHN425_map_data_9);
  FE_PHC424_map_data_21 : CKBD0BWP7T port map(I => map_data(21), Z => FE_PHN424_map_data_21);
  FE_PHC423_map_data_26 : CKBD0BWP7T port map(I => FE_PHN504_map_data_26, Z => FE_PHN423_map_data_26);
  FE_PHC422_map_data_41 : CKBD0BWP7T port map(I => map_data(41), Z => FE_PHN422_map_data_41);
  FE_PHC421_spi_com_MISO_shift_18 : DEL01BWP7T port map(I => FE_PHN421_spi_com_MISO_shift_18, Z => FE_PHN172_spi_com_MISO_shift_18);
  FE_PHC420_spi_com_n_74 : CKBD0BWP7T port map(I => spi_com_n_74, Z => FE_PHN420_spi_com_n_74);
  FE_PHC419_spi_com_bit_count_0 : DEL01BWP7T port map(I => FE_PHN374_spi_com_bit_count_0, Z => FE_PHN419_spi_com_bit_count_0);
  FE_PHC418_spi_com_MISO_shift_46 : DEL01BWP7T port map(I => FE_PHN418_spi_com_MISO_shift_46, Z => FE_PHN368_spi_com_MISO_shift_46);
  FE_PHC417_map_data_8 : CKBD2BWP7T port map(I => FE_PHN390_map_data_8, Z => FE_PHN417_map_data_8);
  FE_PHC416_map_data_58 : BUFFD3BWP7T port map(I => FE_PHN388_map_data_58, Z => FE_PHN416_map_data_58);
  FE_PHC415_map_data_2 : CKBD2BWP7T port map(I => FE_PHN389_map_data_2, Z => FE_PHN415_map_data_2);
  FE_PHC414_map_data_4 : CKBD2BWP7T port map(I => FE_PHN384_map_data_4, Z => FE_PHN414_map_data_4);
  FE_PHC413_level_d_4 : DEL02BWP7T port map(I => FE_PHN382_level_d_4, Z => FE_PHN413_level_d_4);
  FE_PHC412_stable_map_com_n_84 : CKBD0BWP7T port map(I => stable_map_com_n_84, Z => FE_PHN412_stable_map_com_n_84);
  FE_PHC411_map_data_6 : CKBD0BWP7T port map(I => FE_PHN392_map_data_6, Z => FE_PHN411_map_data_6);
  FE_PHC410_energy_d_11 : CKBD2BWP7T port map(I => energy_d(11), Z => FE_PHN410_energy_d_11);
  FE_PHC409_spi_com_MISO_shift_11 : DEL01BWP7T port map(I => spi_com_MISO_shift(11), Z => FE_PHN409_spi_com_MISO_shift_11);
  FE_PHC408_vga_com_texture_module_n_193 : DEL01BWP7T port map(I => vga_com_texture_module_n_193, Z => FE_PHN408_vga_com_texture_module_n_193);
  FE_PHC407_fsm_com_n_106 : DEL02BWP7T port map(I => fsm_com_n_106, Z => FE_PHN407_fsm_com_n_106);
  FE_PHC406_spi_com_n_178 : CKBD2BWP7T port map(I => FE_PHN406_spi_com_n_178, Z => spi_com_n_178);
  FE_PHC405_spi_com_n_83 : CKBD0BWP7T port map(I => spi_com_n_83, Z => FE_PHN405_spi_com_n_83);
  FE_PHC404_vga_com_texture_module_n_252 : DEL0BWP7T port map(I => FE_PHN404_vga_com_texture_module_n_252, Z => vga_com_texture_module_n_252);
  FE_PHC403_energy_d_1 : DEL2BWP7T port map(I => energy_d(1), Z => FE_PHN403_energy_d_1);
  FE_PHC402_energy_d_11 : DEL02BWP7T port map(I => FE_PHN402_energy_d_11, Z => energy_d(11));
  FE_PHC401_vga_com_vcount_2 : CKBD0BWP7T port map(I => FE_PHN401_vga_com_vcount_2, Z => vga_com_vcount(2));
  FE_PHC400_energy_d_7 : CKBD0BWP7T port map(I => energy_d(7), Z => FE_PHN400_energy_d_7);
  FE_PHC399_fsm_com_energy_8 : DEL01BWP7T port map(I => fsm_com_energy(8), Z => FE_PHN399_fsm_com_energy_8);
  FE_PHC398_spi_com_MISO_shift_18 : CKBD2BWP7T port map(I => spi_com_MISO_shift(18), Z => FE_PHN398_spi_com_MISO_shift_18);
  FE_PHC397_fsm_com_energy_0 : DEL01BWP7T port map(I => fsm_com_energy(0), Z => FE_PHN397_fsm_com_energy_0);
  FE_PHC396_fsm_com_reached_high_0 : DEL01BWP7T port map(I => FE_PHN224_fsm_com_reached_high_0, Z => FE_PHN396_fsm_com_reached_high_0);
  FE_PHC395_fsm_com_energy_3 : DEL01BWP7T port map(I => FE_PHN221_fsm_com_energy_3, Z => FE_PHN395_fsm_com_energy_3);
  FE_PHC394_map_data_64 : CKBD0BWP7T port map(I => map_data(64), Z => FE_PHN394_map_data_64);
  FE_PHC393_stable_map_com_n_84 : CKBD0BWP7T port map(I => FE_PHN393_stable_map_com_n_84, Z => stable_map_com_n_84);
  FE_PHC392_map_data_6 : CKBD0BWP7T port map(I => map_data(6), Z => FE_PHN392_map_data_6);
  FE_PHC391_vga_com_texture_module_vvis_0 : DEL01BWP7T port map(I => vga_com_texture_module_vvis(0), Z => FE_PHN391_vga_com_texture_module_vvis_0);
  FE_PHC390_map_data_8 : CKBD2BWP7T port map(I => map_data(8), Z => FE_PHN390_map_data_8);
  FE_PHC389_map_data_2 : CKBD2BWP7T port map(I => map_data(2), Z => FE_PHN389_map_data_2);
  FE_PHC388_map_data_58 : CKBD2BWP7T port map(I => map_data(58), Z => FE_PHN388_map_data_58);
  FE_PHC387_map_data_62 : DEL01BWP7T port map(I => map_data(62), Z => FE_PHN387_map_data_62);
  FE_PHC386_vga_com_texture_module_n_129 : DEL01BWP7T port map(I => FE_PHN220_vga_com_texture_module_n_129, Z => FE_PHN386_vga_com_texture_module_n_129);
  FE_PHC385_map_data_volatile_71 : DEL01BWP7T port map(I => map_data_volatile(71), Z => FE_PHN385_map_data_volatile_71);
  FE_PHC384_map_data_4 : BUFFD0BWP7T port map(I => FE_PHN465_map_data_4, Z => FE_PHN384_map_data_4);
  FE_PHC383_energy_d_10 : CKBD0BWP7T port map(I => energy_d(10), Z => FE_PHN383_energy_d_10);
  FE_PHC382_level_d_4 : BUFFD0BWP7T port map(I => level_d(4), Z => FE_PHN382_level_d_4);
  FE_PHC381_map_data_volatile_46 : DEL01BWP7T port map(I => FE_PHN179_map_data_volatile_46, Z => FE_PHN381_map_data_volatile_46);
  FE_PHC380_spi_com_MISO_shift_40 : DEL01BWP7T port map(I => spi_com_MISO_shift(40), Z => FE_PHN380_spi_com_MISO_shift_40);
  FE_PHC379_spi_com_MOSI_shift_14 : DEL01BWP7T port map(I => FE_PHN379_spi_com_MOSI_shift_14, Z => FE_PHN182_spi_com_MOSI_shift_14);
  FE_PHC378_map_data_volatile_37 : DEL01BWP7T port map(I => FE_PHN181_map_data_volatile_37, Z => FE_PHN378_map_data_volatile_37);
  FE_PHC377_map_data_volatile_36 : DEL01BWP7T port map(I => map_data_volatile(36), Z => FE_PHN377_map_data_volatile_36);
  FE_PHC376_spi_com_MISO_shift_12 : CKBD0BWP7T port map(I => spi_com_MISO_shift(12), Z => FE_PHN376_spi_com_MISO_shift_12);
  FE_PHC375_spi_com_MOSI_shift_12 : DEL01BWP7T port map(I => FE_PHN375_spi_com_MOSI_shift_12, Z => FE_PHN192_spi_com_MOSI_shift_12);
  FE_PHC374_spi_com_bit_count_0 : CKBD0BWP7T port map(I => FE_PHN226_spi_com_bit_count_0, Z => FE_PHN374_spi_com_bit_count_0);
  FE_PHC373_n_87 : DEL01BWP7T port map(I => FE_PHN373_n_87, Z => FE_PHN198_n_87);
  FE_PHC372_n_95 : DEL01BWP7T port map(I => n_95, Z => FE_PHN372_n_95);
  FE_PHC371_spi_com_SCLK_count_1 : BUFFD1P5BWP7T port map(I => FE_PHN240_spi_com_SCLK_count_1, Z => FE_PHN371_spi_com_SCLK_count_1);
  FE_PHC370_vga_com_texture_module_hvis_3 : CKBD3BWP7T port map(I => FE_PHN251_vga_com_texture_module_hvis_3, Z => FE_PHN370_vga_com_texture_module_hvis_3);
  FE_PHC369_spi_com_MISO_shift_34 : CKBD0BWP7T port map(I => FE_PHN369_spi_com_MISO_shift_34, Z => FE_PHN185_spi_com_MISO_shift_34);
  FE_PHC368_spi_com_MISO_shift_46 : CKBD0BWP7T port map(I => FE_PHN368_spi_com_MISO_shift_46, Z => FE_PHN191_spi_com_MISO_shift_46);
  FE_PHC367_spi_com_MISO_shift_14 : CKBD0BWP7T port map(I => spi_com_MISO_shift(14), Z => FE_PHN367_spi_com_MISO_shift_14);
  FE_PHC366_spi_com_MISO_shift_42 : DEL02BWP7T port map(I => FE_PHN366_spi_com_MISO_shift_42, Z => spi_com_MISO_shift(42));
  FE_PHC365_fsm_com_n_20 : CKBD0BWP7T port map(I => FE_PHN365_fsm_com_n_20, Z => fsm_com_n_20);
  FE_PHC364_map_data_volatile_10 : DEL0BWP7T port map(I => FE_PHN364_map_data_volatile_10, Z => map_data_volatile(10));
  FE_PHC363_fsm_com_n_103 : DEL01BWP7T port map(I => fsm_com_n_103, Z => FE_PHN363_fsm_com_n_103);
  FE_PHC362_vga_com_texture_module_n_176 : DEL01BWP7T port map(I => vga_com_texture_module_n_176, Z => FE_PHN362_vga_com_texture_module_n_176);
  FE_PHC361_vga_com_texture_module_n_190 : DEL0BWP7T port map(I => vga_com_texture_module_n_190, Z => FE_PHN361_vga_com_texture_module_n_190);
  FE_PHC360_fsm_com_n_497 : DEL0BWP7T port map(I => fsm_com_n_497, Z => FE_PHN360_fsm_com_n_497);
  FE_PHC359_fsm_com_n_225 : DEL0BWP7T port map(I => fsm_com_n_225, Z => FE_PHN359_fsm_com_n_225);
  FE_PHC358_vga_com_texture_module_n_238 : DEL0BWP7T port map(I => vga_com_texture_module_n_238, Z => FE_PHN358_vga_com_texture_module_n_238);
  FE_PHC357_fsm_com_n_298 : DEL0BWP7T port map(I => fsm_com_n_298, Z => FE_PHN357_fsm_com_n_298);
  FE_PHC356_fsm_com_n_197 : DEL0BWP7T port map(I => FE_PHN356_fsm_com_n_197, Z => fsm_com_n_197);
  FE_PHC355_fsm_com_n_482 : DEL0BWP7T port map(I => fsm_com_n_482, Z => FE_PHN355_fsm_com_n_482);
  FE_PHC354_vga_com_texture_module_n_239 : DEL0BWP7T port map(I => vga_com_texture_module_n_239, Z => FE_PHN354_vga_com_texture_module_n_239);
  FE_PHC353_vga_com_texture_module_n_174 : DEL1BWP7T port map(I => vga_com_texture_module_n_174, Z => FE_PHN353_vga_com_texture_module_n_174);
  FE_PHC352_vga_com_texture_module_n_52 : DEL0BWP7T port map(I => vga_com_texture_module_n_52, Z => FE_PHN352_vga_com_texture_module_n_52);
  FE_PHC351_spi_com_n_254 : CKBD0BWP7T port map(I => spi_com_n_254, Z => FE_PHN351_spi_com_n_254);
  FE_PHC350_stable_map_com_n_106 : DEL0BWP7T port map(I => FE_PHN350_stable_map_com_n_106, Z => stable_map_com_n_106);
  FE_PHC349_stable_map_com_n_130 : DEL0BWP7T port map(I => stable_map_com_n_130, Z => FE_PHN349_stable_map_com_n_130);
  FE_PHC348_stable_map_com_n_134 : DEL0BWP7T port map(I => stable_map_com_n_134, Z => FE_PHN348_stable_map_com_n_134);
  FE_PHC347_stable_map_com_n_59 : DEL0BWP7T port map(I => stable_map_com_n_59, Z => FE_PHN347_stable_map_com_n_59);
  FE_PHC346_stable_map_com_n_107 : DEL0BWP7T port map(I => stable_map_com_n_107, Z => FE_PHN346_stable_map_com_n_107);
  FE_PHC345_stable_map_com_n_82 : DEL0BWP7T port map(I => FE_PHN345_stable_map_com_n_82, Z => stable_map_com_n_82);
  FE_PHC344_vga_com_texture_module_n_240 : DEL0BWP7T port map(I => vga_com_texture_module_n_240, Z => FE_PHN344_vga_com_texture_module_n_240);
  FE_PHC343_vga_com_texture_module_n_232 : DEL0BWP7T port map(I => FE_PHN343_vga_com_texture_module_n_232, Z => vga_com_texture_module_n_232);
  FE_PHC342_vga_com_texture_module_n_254 : DEL0BWP7T port map(I => FE_PHN342_vga_com_texture_module_n_254, Z => vga_com_texture_module_n_254);
  FE_PHC341_vga_com_texture_module_n_216 : DEL0BWP7T port map(I => FE_PHN341_vga_com_texture_module_n_216, Z => vga_com_texture_module_n_216);
  FE_PHC340_fsm_com_n_487 : DEL0BWP7T port map(I => fsm_com_n_487, Z => FE_PHN340_fsm_com_n_487);
  FE_PHC339_vga_com_texture_module_n_249 : DEL0BWP7T port map(I => vga_com_texture_module_n_249, Z => FE_PHN339_vga_com_texture_module_n_249);
  FE_PHC338_stable_map_com_n_49 : DEL0BWP7T port map(I => FE_PHN338_stable_map_com_n_49, Z => stable_map_com_n_49);
  FE_PHC337_fsm_com_n_473 : DEL1BWP7T port map(I => fsm_com_n_473, Z => FE_PHN337_fsm_com_n_473);
  FE_PHC336_fsm_com_n_378 : DEL0BWP7T port map(I => FE_PHN336_fsm_com_n_378, Z => fsm_com_n_378);
  FE_PHC335_vga_com_texture_module_n_251 : DEL0BWP7T port map(I => vga_com_texture_module_n_251, Z => FE_PHN335_vga_com_texture_module_n_251);
  FE_PHC334_spi_com_n_45 : DEL0BWP7T port map(I => spi_com_n_45, Z => FE_PHN334_spi_com_n_45);
  FE_PHC333_n_144 : DEL0BWP7T port map(I => n_144, Z => FE_PHN333_n_144);
  FE_PHC332_stable_map_com_n_55 : DEL2BWP7T port map(I => stable_map_com_n_55, Z => FE_PHN332_stable_map_com_n_55);
  FE_PHC331_vga_com_texture_module_n_162 : DEL0BWP7T port map(I => vga_com_texture_module_n_162, Z => FE_PHN331_vga_com_texture_module_n_162);
  FE_PHC330_fsm_com_n_465 : DEL1BWP7T port map(I => FE_PHN330_fsm_com_n_465, Z => fsm_com_n_465);
  FE_PHC329_fsm_com_n_363 : DEL0BWP7T port map(I => fsm_com_n_363, Z => FE_PHN329_fsm_com_n_363);
  FE_PHC328_stable_map_com_n_136 : DEL1BWP7T port map(I => stable_map_com_n_136, Z => FE_PHN328_stable_map_com_n_136);
  FE_PHC327_vga_com_texture_module_n_253 : DEL0BWP7T port map(I => FE_PHN327_vga_com_texture_module_n_253, Z => vga_com_texture_module_n_253);
  FE_PHC326_vga_com_texture_module_n_48 : DEL0BWP7T port map(I => vga_com_texture_module_n_48, Z => FE_PHN326_vga_com_texture_module_n_48);
  FE_PHC325_vga_com_texture_module_n_229 : DEL0BWP7T port map(I => vga_com_texture_module_n_229, Z => FE_PHN325_vga_com_texture_module_n_229);
  FE_PHC324_spi_com_n_246 : DEL1BWP7T port map(I => spi_com_n_246, Z => FE_PHN324_spi_com_n_246);
  FE_PHC323_stable_map_com_n_133 : DEL1BWP7T port map(I => stable_map_com_n_133, Z => FE_PHN323_stable_map_com_n_133);
  FE_PHC322_spi_com_n_257 : DEL1BWP7T port map(I => spi_com_n_257, Z => FE_PHN322_spi_com_n_257);
  FE_PHC321_fsm_com_n_340 : DEL1BWP7T port map(I => fsm_com_n_340, Z => FE_PHN321_fsm_com_n_340);
  FE_PHC320_fsm_com_n_359 : DEL0BWP7T port map(I => fsm_com_n_359, Z => FE_PHN320_fsm_com_n_359);
  FE_PHC319_spi_com_n_258 : DEL1BWP7T port map(I => spi_com_n_258, Z => FE_PHN319_spi_com_n_258);
  FE_PHC318_vga_com_texture_module_n_248 : DEL1BWP7T port map(I => FE_PHN318_vga_com_texture_module_n_248, Z => vga_com_texture_module_n_248);
  FE_PHC317_fsm_com_n_202 : DEL0BWP7T port map(I => fsm_com_n_202, Z => FE_PHN317_fsm_com_n_202);
  FE_PHC316_fsm_com_n_491 : DEL0BWP7T port map(I => fsm_com_n_491, Z => FE_PHN316_fsm_com_n_491);
  FE_PHC315_spi_com_n_224 : DEL1BWP7T port map(I => spi_com_n_224, Z => FE_PHN315_spi_com_n_224);
  FE_PHC314_fsm_com_n_474 : DEL1BWP7T port map(I => fsm_com_n_474, Z => FE_PHN314_fsm_com_n_474);
  FE_PHC313_fsm_com_n_472 : DEL0BWP7T port map(I => FE_PHN313_fsm_com_n_472, Z => fsm_com_n_472);
  FE_PHC312_vga_com_texture_module_n_242 : DEL0BWP7T port map(I => vga_com_texture_module_n_242, Z => FE_PHN312_vga_com_texture_module_n_242);
  FE_PHC311_vga_com_texture_module_n_201 : DEL0BWP7T port map(I => vga_com_texture_module_n_201, Z => FE_PHN311_vga_com_texture_module_n_201);
  FE_PHC310_stable_map_com_n_126 : DEL1BWP7T port map(I => stable_map_com_n_126, Z => FE_PHN310_stable_map_com_n_126);
  FE_PHC309_vga_com_texture_module_n_187 : DEL1BWP7T port map(I => FE_PHN309_vga_com_texture_module_n_187, Z => vga_com_texture_module_n_187);
  FE_PHC308_fsm_com_n_380 : CKBD0BWP7T port map(I => fsm_com_n_380, Z => FE_PHN308_fsm_com_n_380);
  FE_PHC307_stable_map_com_n_60 : DEL1BWP7T port map(I => stable_map_com_n_60, Z => FE_PHN307_stable_map_com_n_60);
  FE_PHC306_spi_com_n_243 : DEL1BWP7T port map(I => FE_PHN306_spi_com_n_243, Z => spi_com_n_243);
  FE_PHC305_stable_map_com_n_137 : DEL0BWP7T port map(I => stable_map_com_n_137, Z => FE_PHN305_stable_map_com_n_137);
  FE_PHC304_fsm_com_n_477 : DEL1BWP7T port map(I => fsm_com_n_477, Z => FE_PHN304_fsm_com_n_477);
  FE_PHC303_spi_com_n_55 : DEL1BWP7T port map(I => spi_com_n_55, Z => FE_PHN303_spi_com_n_55);
  FE_PHC302_spi_com_n_226 : DEL1BWP7T port map(I => spi_com_n_226, Z => FE_PHN302_spi_com_n_226);
  FE_PHC301_spi_com_n_242 : DEL1BWP7T port map(I => FE_PHN301_spi_com_n_242, Z => spi_com_n_242);
  FE_PHC300_vga_com_texture_module_n_223 : DEL0BWP7T port map(I => FE_PHN300_vga_com_texture_module_n_223, Z => vga_com_texture_module_n_223);
  FE_PHC299_fsm_com_n_357 : DEL0BWP7T port map(I => fsm_com_n_357, Z => FE_PHN299_fsm_com_n_357);
  FE_PHC298_vga_com_texture_module_n_202 : DEL0BWP7T port map(I => vga_com_texture_module_n_202, Z => FE_PHN298_vga_com_texture_module_n_202);
  FE_PHC297_stable_map_com_n_109 : DEL1BWP7T port map(I => stable_map_com_n_109, Z => FE_PHN297_stable_map_com_n_109);
  FE_PHC296_fsm_com_n_464 : DEL0BWP7T port map(I => fsm_com_n_464, Z => FE_PHN296_fsm_com_n_464);
  FE_PHC295_spi_com_n_229 : DEL1BWP7T port map(I => FE_PHN295_spi_com_n_229, Z => spi_com_n_229);
  FE_PHC294_spi_com_n_247 : DEL1BWP7T port map(I => spi_com_n_247, Z => FE_PHN294_spi_com_n_247);
  FE_PHC293_stable_map_com_n_72 : DEL1BWP7T port map(I => stable_map_com_n_72, Z => FE_PHN293_stable_map_com_n_72);
  FE_PHC292_spi_com_n_43 : DEL1BWP7T port map(I => spi_com_n_43, Z => FE_PHN292_spi_com_n_43);
  FE_PHC291_fsm_com_n_485 : DEL0BWP7T port map(I => fsm_com_n_485, Z => FE_PHN291_fsm_com_n_485);
  FE_PHC290_spi_com_n_101 : DEL1BWP7T port map(I => spi_com_n_101, Z => FE_PHN290_spi_com_n_101);
  FE_PHC289_stable_map_com_n_98 : DEL1BWP7T port map(I => stable_map_com_n_98, Z => FE_PHN289_stable_map_com_n_98);
  FE_PHC288_spi_com_n_129 : DEL1BWP7T port map(I => spi_com_n_129, Z => FE_PHN288_spi_com_n_129);
  FE_PHC287_stable_map_com_n_111 : DEL1BWP7T port map(I => stable_map_com_n_111, Z => FE_PHN287_stable_map_com_n_111);
  FE_PHC286_fsm_com_n_429 : DEL0BWP7T port map(I => fsm_com_n_429, Z => FE_PHN286_fsm_com_n_429);
  FE_PHC285_stable_map_com_n_76 : DEL1BWP7T port map(I => stable_map_com_n_76, Z => FE_PHN285_stable_map_com_n_76);
  FE_PHC284_stable_map_com_n_90 : DEL1BWP7T port map(I => FE_PHN284_stable_map_com_n_90, Z => stable_map_com_n_90);
  FE_PHC283_stable_map_com_n_129 : DEL1BWP7T port map(I => FE_PHN283_stable_map_com_n_129, Z => stable_map_com_n_129);
  FE_PHC282_fsm_com_n_466 : DEL0BWP7T port map(I => fsm_com_n_466, Z => FE_PHN282_fsm_com_n_466);
  FE_PHC281_vga_com_texture_module_n_244 : DEL0BWP7T port map(I => vga_com_texture_module_n_244, Z => FE_PHN281_vga_com_texture_module_n_244);
  FE_PHC280_stable_map_com_n_108 : DEL1BWP7T port map(I => stable_map_com_n_108, Z => FE_PHN280_stable_map_com_n_108);
  FE_PHC279_spi_com_n_256 : DEL1BWP7T port map(I => spi_com_n_256, Z => FE_PHN279_spi_com_n_256);
  FE_PHC278_stable_map_com_n_135 : DEL0BWP7T port map(I => stable_map_com_n_135, Z => FE_PHN278_stable_map_com_n_135);
  FE_PHC277_stable_map_com_n_67 : DEL1BWP7T port map(I => FE_PHN277_stable_map_com_n_67, Z => stable_map_com_n_67);
  FE_PHC276_stable_map_com_n_71 : DEL1BWP7T port map(I => stable_map_com_n_71, Z => FE_PHN276_stable_map_com_n_71);
  FE_PHC275_spi_com_n_260 : DEL1BWP7T port map(I => spi_com_n_260, Z => FE_PHN275_spi_com_n_260);
  FE_PHC274_stable_map_com_n_73 : DEL1BWP7T port map(I => stable_map_com_n_73, Z => FE_PHN274_stable_map_com_n_73);
  FE_PHC273_stable_map_com_n_78 : DEL1BWP7T port map(I => FE_PHN273_stable_map_com_n_78, Z => stable_map_com_n_78);
  FE_PHC272_stable_map_com_n_56 : DEL1BWP7T port map(I => stable_map_com_n_56, Z => FE_PHN272_stable_map_com_n_56);
  FE_PHC271_stable_map_com_n_127 : DEL0BWP7T port map(I => stable_map_com_n_127, Z => FE_PHN271_stable_map_com_n_127);
  FE_PHC270_stable_map_com_n_68 : DEL1BWP7T port map(I => FE_PHN270_stable_map_com_n_68, Z => stable_map_com_n_68);
  FE_PHC269_spi_com_n_252 : DEL0BWP7T port map(I => spi_com_n_252, Z => FE_PHN269_spi_com_n_252);
  FE_PHC268_stable_map_com_n_128 : DEL0BWP7T port map(I => FE_PHN268_stable_map_com_n_128, Z => stable_map_com_n_128);
  FE_PHC267_stable_map_com_n_139 : DEL0BWP7T port map(I => FE_PHN267_stable_map_com_n_139, Z => stable_map_com_n_139);
  FE_PHC266_fsm_com_n_337 : DEL0BWP7T port map(I => FE_PHN266_fsm_com_n_337, Z => fsm_com_n_337);
  FE_PHC265_spi_com_n_175 : DEL0BWP7T port map(I => spi_com_n_175, Z => FE_PHN265_spi_com_n_175);
  FE_PHC264_fsm_com_n_483 : DEL0BWP7T port map(I => fsm_com_n_483, Z => FE_PHN264_fsm_com_n_483);
  FE_PHC263_stable_map_com_n_138 : DEL0BWP7T port map(I => FE_PHN263_stable_map_com_n_138, Z => stable_map_com_n_138);
  FE_PHC262_fsm_com_n_434 : DEL0BWP7T port map(I => fsm_com_n_434, Z => FE_PHN262_fsm_com_n_434);
  FE_PHC261_spi_com_n_182 : DEL0BWP7T port map(I => spi_com_n_182, Z => FE_PHN261_spi_com_n_182);
  FE_PHC260_spi_com_n_255 : DEL0BWP7T port map(I => spi_com_n_255, Z => FE_PHN260_spi_com_n_255);
  FE_PHC259_vga_com_texture_module_n_247 : DEL0BWP7T port map(I => vga_com_texture_module_n_247, Z => FE_PHN259_vga_com_texture_module_n_247);
  FE_PHC258_stable_map_com_n_92 : DEL0BWP7T port map(I => stable_map_com_n_92, Z => FE_PHN258_stable_map_com_n_92);
  FE_PHC257_stable_map_com_n_104 : DEL0BWP7T port map(I => stable_map_com_n_104, Z => FE_PHN257_stable_map_com_n_104);
  FE_PHC256_spi_com_n_261 : DEL1BWP7T port map(I => spi_com_n_261, Z => FE_PHN256_spi_com_n_261);
  FE_PHC255_spi_com_n_262 : DEL0BWP7T port map(I => spi_com_n_262, Z => FE_PHN255_spi_com_n_262);
  FE_PHC254_vga_com_texture_module_xposition_4 : DEL02BWP7T port map(I => FE_PHN254_vga_com_texture_module_xposition_4, Z => vga_com_texture_module_xposition(4));
  FE_PHC253_vga_com_texture_module_yposition_0 : DEL01BWP7T port map(I => vga_com_texture_module_yposition(0), Z => FE_PHN253_vga_com_texture_module_yposition_0);
  FE_PHC252_vga_com_texture_module_vvis_0 : DEL02BWP7T port map(I => FE_PHN252_vga_com_texture_module_vvis_0, Z => vga_com_texture_module_vvis(0));
  FE_PHC251_vga_com_texture_module_hvis_3 : DEL02BWP7T port map(I => vga_com_texture_module_hvis(3), Z => FE_PHN251_vga_com_texture_module_hvis_3);
  FE_PHC250_level_d_0 : DEL0BWP7T port map(I => FE_PHN250_level_d_0, Z => level_d(0));
  FE_PHC249_score_d_8 : DEL1BWP7T port map(I => score_d(8), Z => FE_PHN249_score_d_8);
  FE_PHC248_energy_d_4 : DEL0BWP7T port map(I => FE_PHN248_energy_d_4, Z => energy_d(4));
  FE_PHC247_energy_d_0 : DEL0BWP7T port map(I => FE_PHN247_energy_d_0, Z => energy_d(0));
  FE_PHC246_energy_d_1 : DEL02BWP7T port map(I => FE_PHN246_energy_d_1, Z => energy_d(1));
  FE_PHC245_energy_d_8 : DEL0BWP7T port map(I => FE_PHN245_energy_d_8, Z => energy_d(8));
  FE_PHC244_score_d_4 : DEL0BWP7T port map(I => score_d(4), Z => FE_PHN244_score_d_4);
  FE_PHC243_level_abs_0 : DEL02BWP7T port map(I => FE_PHN243_level_abs_0, Z => level_abs(0));
  FE_PHC242_vga_com_vcount_5 : DEL2BWP7T port map(I => FE_PHN242_vga_com_vcount_5, Z => vga_com_vcount(5));
  FE_PHC241_vga_com_vcount_9 : DEL1BWP7T port map(I => vga_com_vcount(9), Z => FE_PHN241_vga_com_vcount_9);
  FE_PHC240_spi_com_SCLK_count_1 : CKBD0BWP7T port map(I => spi_com_SCLK_count(1), Z => FE_PHN240_spi_com_SCLK_count_1);
  FE_PHC239_vga_com_vcount_8 : DEL1BWP7T port map(I => vga_com_vcount(8), Z => FE_PHN239_vga_com_vcount_8);
  FE_PHC238_vga_com_vcount_7 : DEL0BWP7T port map(I => vga_com_vcount(7), Z => FE_PHN238_vga_com_vcount_7);
  FE_PHC237_spi_com_state_2 : DEL02BWP7T port map(I => spi_com_state(2), Z => FE_PHN237_spi_com_state_2);
  FE_PHC236_vga_com_hcount_8 : DEL02BWP7T port map(I => FE_PHN236_vga_com_hcount_8, Z => vga_com_hcount(8));
  FE_PHC235_vga_com_hcount_9 : DEL02BWP7T port map(I => vga_com_hcount(9), Z => FE_PHN235_vga_com_hcount_9);
  FE_PHC234_vga_com_vcount_6 : DEL1BWP7T port map(I => FE_PHN234_vga_com_vcount_6, Z => vga_com_vcount(6));
  FE_PHC233_fsm_com_n_22 : DEL01BWP7T port map(I => fsm_com_n_22, Z => FE_PHN233_fsm_com_n_22);
  FE_PHC232_energy_d_7 : DEL02BWP7T port map(I => FE_PHN400_energy_d_7, Z => FE_PHN232_energy_d_7);
  FE_PHC231_vga_com_vcount_2 : DEL02BWP7T port map(I => vga_com_vcount(2), Z => FE_PHN231_vga_com_vcount_2);
  FE_PHC230_fsm_com_energy_2 : DEL01BWP7T port map(I => fsm_com_energy(2), Z => FE_PHN230_fsm_com_energy_2);
  FE_PHC229_spi_com_SCLK_count_0 : DEL1BWP7T port map(I => spi_com_SCLK_count(0), Z => FE_PHN229_spi_com_SCLK_count_0);
  FE_PHC228_spi_com_byte_count_0 : DEL1BWP7T port map(I => FE_PHN228_spi_com_byte_count_0, Z => spi_com_byte_count(0));
  FE_PHC227_score_d_12 : DEL1BWP7T port map(I => score_d(12), Z => FE_PHN227_score_d_12);
  FE_PHC226_spi_com_bit_count_0 : DEL02BWP7T port map(I => spi_com_bit_count(0), Z => FE_PHN226_spi_com_bit_count_0);
  FE_PHC225_fsm_com_energy_8 : CKBD0BWP7T port map(I => FE_PHN399_fsm_com_energy_8, Z => FE_PHN225_fsm_com_energy_8);
  FE_PHC224_fsm_com_reached_high_0 : DEL02BWP7T port map(I => fsm_com_reached_high(0), Z => FE_PHN224_fsm_com_reached_high_0);
  FE_PHC223_fsm_com_n_8 : DEL01BWP7T port map(I => fsm_com_n_8, Z => FE_PHN223_fsm_com_n_8);
  FE_PHC222_vga_com_display_controller_module_display_state_0 : DEL01BWP7T port map(I => vga_com_display_controller_module_display_state(0), Z => FE_PHN222_vga_com_display_controller_module_display_state_0);
  FE_PHC221_fsm_com_energy_3 : CKBD0BWP7T port map(I => fsm_com_energy(3), Z => FE_PHN221_fsm_com_energy_3);
  FE_PHC220_vga_com_texture_module_n_129 : CKBD0BWP7T port map(I => vga_com_texture_module_n_129, Z => FE_PHN220_vga_com_texture_module_n_129);
  FE_PHC219_vga_com_texture_module_n_134 : DEL0BWP7T port map(I => FE_PHN219_vga_com_texture_module_n_134, Z => vga_com_texture_module_n_134);
  FE_PHC218_spi_com_pause_count_0 : DEL1BWP7T port map(I => FE_PHN218_spi_com_pause_count_0, Z => spi_com_pause_count(0));
  FE_PHC217_vga_com_texture_module_n_6 : DEL1BWP7T port map(I => vga_com_texture_module_n_6, Z => FE_PHN217_vga_com_texture_module_n_6);
  FE_PHC216_vga_com_texture_module_n_115 : CKBD3BWP7T port map(I => vga_com_texture_module_n_115, Z => FE_PHN216_vga_com_texture_module_n_115);
  FE_PHC215_fsm_com_n_6 : DEL0BWP7T port map(I => fsm_com_n_6, Z => FE_PHN215_fsm_com_n_6);
  FE_PHC214_energy_d_3 : DEL0BWP7T port map(I => energy_d(3), Z => FE_PHN214_energy_d_3);
  FE_PHC213_vga_com_texture_module_n_204 : DEL0BWP7T port map(I => vga_com_texture_module_n_204, Z => FE_PHN213_vga_com_texture_module_n_204);
  FE_PHC212_fsm_com_edge_detec2_3 : DEL1BWP7T port map(I => fsm_com_edge_detec2(3), Z => FE_PHN212_fsm_com_edge_detec2_3);
  FE_PHC211_vga_com_hcount_6 : CKBD0BWP7T port map(I => vga_com_hcount(6), Z => FE_PHN211_vga_com_hcount_6);
  FE_PHC210_fsm_com_edge_detec1_3 : DEL1BWP7T port map(I => FE_PHN210_fsm_com_edge_detec1_3, Z => fsm_com_edge_detec1(3));
  FE_PHC209_fsm_com_edge_detec0_3 : DEL1BWP7T port map(I => fsm_com_edge_detec0(3), Z => FE_PHN209_fsm_com_edge_detec0_3);
  FE_PHC208_fsm_com_n_20 : DEL02BWP7T port map(I => fsm_com_n_20, Z => FE_PHN208_fsm_com_n_20);
  FE_PHC207_button_left : DEL0BWP7T port map(I => button_left, Z => FE_PHN207_button_left);
  FE_PHC206_fsm_com_energy_7 : DEL0BWP7T port map(I => fsm_com_energy(7), Z => FE_PHN206_fsm_com_energy_7);
  FE_PHC205_fsm_com_reached_high_1 : DEL02BWP7T port map(I => fsm_com_reached_high(1), Z => FE_PHN205_fsm_com_reached_high_1);
  FE_PHC204_vga_com_texture_module_n_16 : DEL0BWP7T port map(I => FE_PHN204_vga_com_texture_module_n_16, Z => vga_com_texture_module_n_16);
  FE_PHC203_vga_com_texture_module_n_79 : DEL0BWP7T port map(I => vga_com_texture_module_n_79, Z => FE_PHN203_vga_com_texture_module_n_79);
  FE_PHC202_fsm_com_energy_4 : DEL0BWP7T port map(I => fsm_com_energy(4), Z => FE_PHN202_fsm_com_energy_4);
  FE_PHC201_n_95 : DEL0BWP7T port map(I => FE_PHN372_n_95, Z => FE_PHN201_n_95);
  FE_PHC200_vga_com_vcount_0 : DEL1BWP7T port map(I => vga_com_vcount(0), Z => FE_PHN200_vga_com_vcount_0);
  FE_PHC199_vga_com_texture_module_n_18 : DEL0BWP7T port map(I => vga_com_texture_module_n_18, Z => FE_PHN199_vga_com_texture_module_n_18);
  FE_PHC198_n_87 : DEL0BWP7T port map(I => FE_PHN198_n_87, Z => n_87);
  FE_PHC197_vga_com_texture_module_n_105 : DEL0BWP7T port map(I => FE_PHN197_vga_com_texture_module_n_105, Z => vga_com_texture_module_n_105);
  FE_PHC196_button_right : DEL0BWP7T port map(I => button_right, Z => FE_PHN196_button_right);
  FE_PHC195_button_up : DEL0BWP7T port map(I => button_up, Z => FE_PHN195_button_up);
  FE_PHC194_vga_com_texture_module_n_164 : DEL0BWP7T port map(I => vga_com_texture_module_n_164, Z => FE_PHN194_vga_com_texture_module_n_164);
  FE_PHC193_vga_com_texture_module_n_17 : DEL1BWP7T port map(I => vga_com_texture_module_n_17, Z => FE_PHN193_vga_com_texture_module_n_17);
  FE_PHC192_spi_com_MOSI_shift_12 : DEL02BWP7T port map(I => FE_PHN192_spi_com_MOSI_shift_12, Z => spi_com_MOSI_shift(12));
  FE_PHC191_spi_com_MISO_shift_46 : DEL02BWP7T port map(I => FE_PHN191_spi_com_MISO_shift_46, Z => spi_com_MISO_shift(46));
  FE_PHC190_spi_com_MISO_shift_14 : DEL02BWP7T port map(I => FE_PHN367_spi_com_MISO_shift_14, Z => FE_PHN190_spi_com_MISO_shift_14);
  FE_PHC189_energy_d_2 : DEL0BWP7T port map(I => energy_d(2), Z => FE_PHN189_energy_d_2);
  FE_PHC188_fsm_com_n_28 : DEL1BWP7T port map(I => fsm_com_n_28, Z => FE_PHN188_fsm_com_n_28);
  FE_PHC187_spi_com_MISO_shift_12 : DEL02BWP7T port map(I => FE_PHN376_spi_com_MISO_shift_12, Z => FE_PHN187_spi_com_MISO_shift_12);
  FE_PHC186_n_93 : DEL2BWP7T port map(I => n_93, Z => FE_PHN186_n_93);
  FE_PHC185_spi_com_MISO_shift_34 : DEL02BWP7T port map(I => FE_PHN185_spi_com_MISO_shift_34, Z => spi_com_MISO_shift(34));
  FE_PHC184_fsm_com_n_27 : DEL1BWP7T port map(I => fsm_com_n_27, Z => FE_PHN184_fsm_com_n_27);
  FE_PHC183_map_data_volatile_33 : DEL0BWP7T port map(I => FE_PHN183_map_data_volatile_33, Z => map_data_volatile(33));
  FE_PHC182_spi_com_MOSI_shift_14 : DEL0BWP7T port map(I => FE_PHN182_spi_com_MOSI_shift_14, Z => spi_com_MOSI_shift(14));
  FE_PHC181_map_data_volatile_37 : DEL0BWP7T port map(I => map_data_volatile(37), Z => FE_PHN181_map_data_volatile_37);
  FE_PHC180_spi_com_n_5 : DEL1BWP7T port map(I => FE_PHN180_spi_com_n_5, Z => spi_com_n_5);
  FE_PHC179_map_data_volatile_46 : DEL0BWP7T port map(I => map_data_volatile(46), Z => FE_PHN179_map_data_volatile_46);
  FE_PHC178_map_data_volatile_36 : DEL0BWP7T port map(I => FE_PHN178_map_data_volatile_36, Z => map_data_volatile(36));
  FE_PHC177_map_data_volatile_71 : DEL0BWP7T port map(I => FE_PHN177_map_data_volatile_71, Z => map_data_volatile(71));
  FE_PHC176_stable_map_com_n_35 : DEL0BWP7T port map(I => stable_map_com_n_35, Z => FE_PHN176_stable_map_com_n_35);
  FE_PHC175_spi_com_n_9 : DEL1BWP7T port map(I => spi_com_n_9, Z => FE_PHN175_spi_com_n_9);
  FE_PHC174_score_d_1 : DEL0BWP7T port map(I => score_d(1), Z => FE_PHN174_score_d_1);
  FE_PHC173_spi_com_MISO_shift_11 : DEL02BWP7T port map(I => FE_PHN173_spi_com_MISO_shift_11, Z => spi_com_MISO_shift(11));
  FE_PHC172_spi_com_MISO_shift_18 : DEL02BWP7T port map(I => FE_PHN172_spi_com_MISO_shift_18, Z => spi_com_MISO_shift(18));
  FE_PHC171_map_data_10 : DEL1BWP7T port map(I => map_data(10), Z => FE_PHN171_map_data_10);
  FE_PHC170_spi_com_MISO_shift_40 : DEL0BWP7T port map(I => FE_PHN380_spi_com_MISO_shift_40, Z => FE_PHN170_spi_com_MISO_shift_40);
  FE_PHC169_n_86 : DEL1BWP7T port map(I => n_86, Z => FE_PHN169_n_86);
  FE_PHC168_n_91 : DEL1BWP7T port map(I => n_91, Z => FE_PHN168_n_91);
  FE_PHC167_n_94 : DEL1BWP7T port map(I => FE_PHN167_n_94, Z => n_94);
  FE_PHC166_n_90 : DEL1BWP7T port map(I => n_90, Z => FE_PHN166_n_90);
  FE_PHC165_n_96 : DEL1BWP7T port map(I => FE_PHN165_n_96, Z => n_96);
  FE_PHC164_n_92 : DEL1BWP7T port map(I => FE_PHN164_n_92, Z => n_92);
  FE_PHC163_n_85 : DEL1BWP7T port map(I => FE_PHN163_n_85, Z => n_85);
  FE_PHC162_spi_com_MISO_shift_3 : DEL2BWP7T port map(I => FE_PHN162_spi_com_MISO_shift_3, Z => spi_com_MISO_shift(3));
  FE_PHC161_vga_com_hcount_7 : DEL02BWP7T port map(I => vga_com_hcount(7), Z => FE_PHN161_vga_com_hcount_7);
  FE_PHC160_n_89 : DEL1BWP7T port map(I => n_89, Z => FE_PHN160_n_89);
  FE_PHC159_n_88 : DEL1BWP7T port map(I => FE_PHN159_n_88, Z => n_88);
  FE_PHC158_map_data_volatile_58 : DEL2BWP7T port map(I => FE_PHN158_map_data_volatile_58, Z => map_data_volatile(58));
  FE_PHC157_map_data_volatile_4 : DEL2BWP7T port map(I => FE_PHN157_map_data_volatile_4, Z => map_data_volatile(4));
  FE_PHC156_spi_com_MISO_shift_49 : DEL2BWP7T port map(I => FE_PHN156_spi_com_MISO_shift_49, Z => spi_com_MISO_shift(49));
  FE_PHC155_spi_com_MISO_shift_44 : DEL2BWP7T port map(I => FE_PHN155_spi_com_MISO_shift_44, Z => spi_com_MISO_shift(44));
  FE_PHC154_map_data_volatile_52 : DEL1BWP7T port map(I => FE_PHN154_map_data_volatile_52, Z => map_data_volatile(52));
  FE_PHC153_spi_com_MISO_shift_47 : DEL1BWP7T port map(I => FE_PHN153_spi_com_MISO_shift_47, Z => spi_com_MISO_shift(47));
  FE_PHC152_spi_com_MISO_shift_39 : DEL1BWP7T port map(I => FE_PHN152_spi_com_MISO_shift_39, Z => spi_com_MISO_shift(39));
  FE_PHC151_spi_com_MISO_shift_64 : DEL0BWP7T port map(I => spi_com_MISO_shift(64), Z => FE_PHN151_spi_com_MISO_shift_64);
  FE_PHC150_map_data_volatile_23 : DEL1BWP7T port map(I => FE_PHN150_map_data_volatile_23, Z => map_data_volatile(23));
  FE_PHC149_spi_com_MISO_shift_62 : DEL1BWP7T port map(I => spi_com_MISO_shift(62), Z => FE_PHN149_spi_com_MISO_shift_62);
  FE_PHC148_spi_com_MISO_shift_51 : DEL0BWP7T port map(I => FE_PHN148_spi_com_MISO_shift_51, Z => spi_com_MISO_shift(51));
  FE_PHC147_map_data_volatile_35 : DEL1BWP7T port map(I => FE_PHN147_map_data_volatile_35, Z => map_data_volatile(35));
  FE_PHC146_spi_com_MOSI_shift_5 : DEL1BWP7T port map(I => FE_PHN146_spi_com_MOSI_shift_5, Z => spi_com_MOSI_shift(5));
  FE_PHC145_spi_com_MISO_shift_27 : DEL1BWP7T port map(I => FE_PHN145_spi_com_MISO_shift_27, Z => spi_com_MISO_shift(27));
  FE_PHC144_spi_com_MISO_shift_0 : DEL1BWP7T port map(I => FE_PHN144_spi_com_MISO_shift_0, Z => spi_com_MISO_shift(0));
  FE_PHC143_fsm_com_n_12 : DEL1BWP7T port map(I => FE_PHN143_fsm_com_n_12, Z => fsm_com_n_12);
  FE_PHC142_spi_com_MOSI_shift_1 : DEL1BWP7T port map(I => FE_PHN142_spi_com_MOSI_shift_1, Z => spi_com_MOSI_shift(1));
  FE_PHC141_spi_com_MOSI_shift_13 : DEL1BWP7T port map(I => spi_com_MOSI_shift(13), Z => FE_PHN141_spi_com_MOSI_shift_13);
  FE_PHC140_spi_com_MISO_shift_13 : DEL1BWP7T port map(I => FE_PHN140_spi_com_MISO_shift_13, Z => spi_com_MISO_shift(13));
  FE_PHC139_map_data_volatile_53 : DEL1BWP7T port map(I => FE_PHN139_map_data_volatile_53, Z => map_data_volatile(53));
  FE_PHC138_spi_com_MISO_shift_33 : DEL0BWP7T port map(I => FE_PHN138_spi_com_MISO_shift_33, Z => spi_com_MISO_shift(33));
  FE_PHC137_map_data_volatile_16 : DEL1BWP7T port map(I => FE_PHN137_map_data_volatile_16, Z => map_data_volatile(16));
  FE_PHC136_fsm_com_edge_detec1_2 : DEL1BWP7T port map(I => fsm_com_edge_detec1(2), Z => FE_PHN136_fsm_com_edge_detec1_2);
  FE_PHC135_spi_com_MISO_shift_1 : DEL0BWP7T port map(I => FE_PHN135_spi_com_MISO_shift_1, Z => spi_com_MISO_shift(1));
  FE_PHC134_map_data_volatile_20 : DEL1BWP7T port map(I => FE_PHN134_map_data_volatile_20, Z => map_data_volatile(20));
  FE_PHC133_map_data_volatile_25 : DEL1BWP7T port map(I => FE_PHN133_map_data_volatile_25, Z => map_data_volatile(25));
  FE_PHC132_map_data_volatile_57 : DEL1BWP7T port map(I => FE_PHN132_map_data_volatile_57, Z => map_data_volatile(57));
  FE_PHC131_spi_com_MOSI_shift_7 : DEL1BWP7T port map(I => FE_PHN131_spi_com_MOSI_shift_7, Z => spi_com_MOSI_shift(7));
  FE_PHC130_map_data_volatile_38 : DEL1BWP7T port map(I => FE_PHN130_map_data_volatile_38, Z => map_data_volatile(38));
  FE_PHC129_spi_com_MOSI_shift_10 : DEL1BWP7T port map(I => FE_PHN129_spi_com_MOSI_shift_10, Z => spi_com_MOSI_shift(10));
  FE_PHC128_spi_com_MOSI_shift_0 : DEL1BWP7T port map(I => FE_PHN128_spi_com_MOSI_shift_0, Z => spi_com_MOSI_shift(0));
  FE_PHC127_map_data_volatile_3 : DEL1BWP7T port map(I => FE_PHN127_map_data_volatile_3, Z => map_data_volatile(3));
  FE_PHC126_map_data_volatile_56 : DEL1BWP7T port map(I => map_data_volatile(56), Z => FE_PHN126_map_data_volatile_56);
  FE_PHC125_map_data_volatile_11 : DEL1BWP7T port map(I => FE_PHN125_map_data_volatile_11, Z => map_data_volatile(11));
  FE_PHC124_map_data_volatile_8 : DEL1BWP7T port map(I => FE_PHN124_map_data_volatile_8, Z => map_data_volatile(8));
  FE_PHC123_fsm_com_edge_detec2_1 : DEL1BWP7T port map(I => fsm_com_edge_detec2(1), Z => FE_PHN123_fsm_com_edge_detec2_1);
  FE_PHC122_map_data_volatile_41 : DEL1BWP7T port map(I => map_data_volatile(41), Z => FE_PHN122_map_data_volatile_41);
  FE_PHC121_spi_com_MISO_shift_17 : DEL1BWP7T port map(I => FE_PHN121_spi_com_MISO_shift_17, Z => spi_com_MISO_shift(17));
  FE_PHC120_fsm_com_edge_detec1_1 : DEL1BWP7T port map(I => fsm_com_edge_detec1(1), Z => FE_PHN120_fsm_com_edge_detec1_1);
  FE_PHC119_map_data_volatile_39 : DEL1BWP7T port map(I => FE_PHN119_map_data_volatile_39, Z => map_data_volatile(39));
  FE_PHC118_map_data_volatile_45 : DEL1BWP7T port map(I => FE_PHN118_map_data_volatile_45, Z => map_data_volatile(45));
  FE_PHC117_spi_com_MISO_shift_52 : DEL1BWP7T port map(I => spi_com_MISO_shift(52), Z => FE_PHN117_spi_com_MISO_shift_52);
  FE_PHC116_map_data_volatile_9 : DEL1BWP7T port map(I => FE_PHN116_map_data_volatile_9, Z => map_data_volatile(9));
  FE_PHC115_spi_com_MISO_shift_61 : DEL1BWP7T port map(I => FE_PHN115_spi_com_MISO_shift_61, Z => spi_com_MISO_shift(61));
  FE_PHC114_spi_com_MISO_shift_50 : DEL1BWP7T port map(I => FE_PHN114_spi_com_MISO_shift_50, Z => spi_com_MISO_shift(50));
  FE_PHC113_map_data_volatile_62 : DEL1BWP7T port map(I => FE_PHN113_map_data_volatile_62, Z => map_data_volatile(62));
  FE_PHC112_spi_com_MOSI_shift_6 : DEL1BWP7T port map(I => spi_com_MOSI_shift(6), Z => FE_PHN112_spi_com_MOSI_shift_6);
  FE_PHC111_map_data_volatile_21 : DEL1BWP7T port map(I => FE_PHN111_map_data_volatile_21, Z => map_data_volatile(21));
  FE_PHC110_map_data_volatile_22 : DEL1BWP7T port map(I => FE_PHN110_map_data_volatile_22, Z => map_data_volatile(22));
  FE_PHC109_map_data_volatile_40 : DEL1BWP7T port map(I => FE_PHN109_map_data_volatile_40, Z => map_data_volatile(40));
  FE_PHC108_map_data_volatile_43 : DEL1BWP7T port map(I => FE_PHN108_map_data_volatile_43, Z => map_data_volatile(43));
  FE_PHC107_spi_com_MISO_shift_57 : DEL1BWP7T port map(I => spi_com_MISO_shift(57), Z => FE_PHN107_spi_com_MISO_shift_57);
  FE_PHC106_map_data_volatile_32 : DEL1BWP7T port map(I => FE_PHN106_map_data_volatile_32, Z => map_data_volatile(32));
  FE_PHC105_fsm_com_edge_detec0_0 : DEL1BWP7T port map(I => fsm_com_edge_detec0(0), Z => FE_PHN105_fsm_com_edge_detec0_0);
  FE_PHC104_map_data_volatile_61 : DEL1BWP7T port map(I => FE_PHN104_map_data_volatile_61, Z => map_data_volatile(61));
  FE_PHC103_spi_com_MISO_shift_58 : DEL1BWP7T port map(I => FE_PHN103_spi_com_MISO_shift_58, Z => spi_com_MISO_shift(58));
  FE_PHC102_spi_com_MISO_shift_65 : DEL1BWP7T port map(I => FE_PHN102_spi_com_MISO_shift_65, Z => spi_com_MISO_shift(65));
  FE_PHC101_vga_com_texture_module_vvis_6 : DEL1BWP7T port map(I => vga_com_texture_module_vvis(6), Z => FE_PHN101_vga_com_texture_module_vvis_6);
  FE_PHC100_fsm_com_edge_detec2_0 : DEL1BWP7T port map(I => fsm_com_edge_detec2(0), Z => FE_PHN100_fsm_com_edge_detec2_0);
  FE_PHC99_map_data_volatile_55 : DEL1BWP7T port map(I => FE_PHN99_map_data_volatile_55, Z => map_data_volatile(55));
  FE_PHC98_map_data_volatile_12 : DEL1BWP7T port map(I => FE_PHN98_map_data_volatile_12, Z => map_data_volatile(12));
  FE_PHC97_spi_com_MISO_shift_9 : DEL1BWP7T port map(I => FE_PHN97_spi_com_MISO_shift_9, Z => spi_com_MISO_shift(9));
  FE_PHC96_spi_com_MOSI_shift_4 : DEL1BWP7T port map(I => spi_com_MOSI_shift(4), Z => FE_PHN96_spi_com_MOSI_shift_4);
  FE_PHC95_map_data_volatile_0 : DEL1BWP7T port map(I => map_data_volatile(0), Z => FE_PHN95_map_data_volatile_0);
  FE_PHC94_map_data_volatile_6 : DEL1BWP7T port map(I => map_data_volatile(6), Z => FE_PHN94_map_data_volatile_6);
  FE_PHC93_fsm_com_edge_detec2_2 : DEL1BWP7T port map(I => fsm_com_edge_detec2(2), Z => FE_PHN93_fsm_com_edge_detec2_2);
  FE_PHC92_spi_com_MOSI_shift_3 : DEL1BWP7T port map(I => spi_com_MOSI_shift(3), Z => FE_PHN92_spi_com_MOSI_shift_3);
  FE_PHC91_fsm_com_edge_detec1_0 : DEL1BWP7T port map(I => fsm_com_edge_detec1(0), Z => FE_PHN91_fsm_com_edge_detec1_0);
  FE_PHC90_map_data_volatile_1 : DEL1BWP7T port map(I => FE_PHN90_map_data_volatile_1, Z => map_data_volatile(1));
  FE_PHC89_map_data_volatile_42 : DEL1BWP7T port map(I => FE_PHN89_map_data_volatile_42, Z => map_data_volatile(42));
  FE_PHC88_map_data_volatile_69 : DEL1BWP7T port map(I => FE_PHN88_map_data_volatile_69, Z => map_data_volatile(69));
  FE_PHC87_spi_com_MISO_shift_55 : DEL1BWP7T port map(I => FE_PHN87_spi_com_MISO_shift_55, Z => spi_com_MISO_shift(55));
  FE_PHC86_map_data_volatile_15 : DEL1BWP7T port map(I => FE_PHN86_map_data_volatile_15, Z => map_data_volatile(15));
  FE_PHC85_map_data_volatile_63 : DEL1BWP7T port map(I => FE_PHN85_map_data_volatile_63, Z => map_data_volatile(63));
  FE_PHC84_map_data_volatile_54 : DEL1BWP7T port map(I => map_data_volatile(54), Z => FE_PHN84_map_data_volatile_54);
  FE_PHC83_spi_com_MISO_shift_28 : DEL0BWP7T port map(I => FE_PHN83_spi_com_MISO_shift_28, Z => spi_com_MISO_shift(28));
  FE_PHC82_map_data_volatile_30 : DEL1BWP7T port map(I => FE_PHN82_map_data_volatile_30, Z => map_data_volatile(30));
  FE_PHC81_spi_com_MISO_shift_72 : DEL1BWP7T port map(I => FE_PHN81_spi_com_MISO_shift_72, Z => spi_com_MISO_shift(72));
  FE_PHC80_fsm_com_edge_detec0_2 : DEL1BWP7T port map(I => fsm_com_edge_detec0(2), Z => FE_PHN80_fsm_com_edge_detec0_2);
  FE_PHC79_fsm_com_edge_detec0_1 : DEL1BWP7T port map(I => fsm_com_edge_detec0(1), Z => FE_PHN79_fsm_com_edge_detec0_1);
  FE_PHC78_map_data_volatile_31 : DEL1BWP7T port map(I => FE_PHN78_map_data_volatile_31, Z => map_data_volatile(31));
  FE_PHC77_map_data_volatile_18 : DEL1BWP7T port map(I => FE_PHN77_map_data_volatile_18, Z => map_data_volatile(18));
  FE_PHC76_map_data_volatile_49 : DEL1BWP7T port map(I => FE_PHN76_map_data_volatile_49, Z => map_data_volatile(49));
  FE_PHC75_spi_com_MOSI_shift_2 : DEL1BWP7T port map(I => spi_com_MOSI_shift(2), Z => FE_PHN75_spi_com_MOSI_shift_2);
  FE_PHC74_map_data_volatile_24 : DEL1BWP7T port map(I => map_data_volatile(24), Z => FE_PHN74_map_data_volatile_24);
  FE_PHC73_map_data_volatile_47 : DEL1BWP7T port map(I => FE_PHN73_map_data_volatile_47, Z => map_data_volatile(47));
  FE_PHC72_spi_com_MISO_shift_20 : DEL1BWP7T port map(I => FE_PHN72_spi_com_MISO_shift_20, Z => spi_com_MISO_shift(20));
  FE_PHC71_map_data_volatile_5 : DEL1BWP7T port map(I => FE_PHN71_map_data_volatile_5, Z => map_data_volatile(5));
  FE_PHC70_map_data_volatile_66 : DEL1BWP7T port map(I => map_data_volatile(66), Z => FE_PHN70_map_data_volatile_66);
  FE_PHC69_spi_com_MISO_shift_25 : DEL1BWP7T port map(I => spi_com_MISO_shift(25), Z => FE_PHN69_spi_com_MISO_shift_25);
  FE_PHC68_spi_com_MISO_shift_10 : DEL1BWP7T port map(I => FE_PHN68_spi_com_MISO_shift_10, Z => spi_com_MISO_shift(10));
  FE_PHC67_spi_com_MISO_shift_45 : DEL1BWP7T port map(I => spi_com_MISO_shift(45), Z => FE_PHN67_spi_com_MISO_shift_45);
  FE_PHC66_spi_com_send_in0 : DEL1BWP7T port map(I => spi_com_send_in0, Z => FE_PHN66_spi_com_send_in0);
  FE_PHC65_map_data_volatile_50 : DEL1BWP7T port map(I => FE_PHN65_map_data_volatile_50, Z => map_data_volatile(50));
  FE_PHC64_spi_com_MISO_shift_6 : DEL1BWP7T port map(I => FE_PHN64_spi_com_MISO_shift_6, Z => spi_com_MISO_shift(6));
  FE_PHC63_map_data_volatile_26 : DEL1BWP7T port map(I => map_data_volatile(26), Z => FE_PHN63_map_data_volatile_26);
  FE_PHC62_spi_com_MISO_shift_32 : DEL1BWP7T port map(I => spi_com_MISO_shift(32), Z => FE_PHN62_spi_com_MISO_shift_32);
  FE_PHC61_map_data_volatile_17 : DEL1BWP7T port map(I => map_data_volatile(17), Z => FE_PHN61_map_data_volatile_17);
  FE_PHC60_map_data_volatile_67 : DEL1BWP7T port map(I => map_data_volatile(67), Z => FE_PHN60_map_data_volatile_67);
  FE_PHC59_map_data_volatile_29 : DEL1BWP7T port map(I => FE_PHN59_map_data_volatile_29, Z => map_data_volatile(29));
  FE_PHC58_map_data_volatile_70 : DEL1BWP7T port map(I => FE_PHN58_map_data_volatile_70, Z => map_data_volatile(70));
  FE_PHC57_spi_com_MISO_shift_35 : DEL1BWP7T port map(I => spi_com_MISO_shift(35), Z => FE_PHN57_spi_com_MISO_shift_35);
  FE_PHC56_map_data_volatile_34 : DEL1BWP7T port map(I => FE_PHN56_map_data_volatile_34, Z => map_data_volatile(34));
  FE_PHC55_map_data_volatile_14 : DEL1BWP7T port map(I => FE_PHN55_map_data_volatile_14, Z => map_data_volatile(14));
  FE_PHC54_spi_com_MISO_shift_43 : DEL1BWP7T port map(I => spi_com_MISO_shift(43), Z => FE_PHN54_spi_com_MISO_shift_43);
  FE_PHC53_spi_com_MISO_shift_26 : DEL1BWP7T port map(I => FE_PHN53_spi_com_MISO_shift_26, Z => spi_com_MISO_shift(26));
  FE_PHC52_map_data_volatile_7 : DEL1BWP7T port map(I => map_data_volatile(7), Z => FE_PHN52_map_data_volatile_7);
  FE_PHC51_spi_com_MISO_shift_41 : DEL1BWP7T port map(I => spi_com_MISO_shift(41), Z => FE_PHN51_spi_com_MISO_shift_41);
  FE_PHC50_map_data_volatile_48 : DEL1BWP7T port map(I => FE_PHN50_map_data_volatile_48, Z => map_data_volatile(48));
  FE_PHC49_map_data_volatile_2 : DEL1BWP7T port map(I => FE_PHN49_map_data_volatile_2, Z => map_data_volatile(2));
  FE_PHC48_map_data_volatile_68 : DEL1BWP7T port map(I => FE_PHN48_map_data_volatile_68, Z => map_data_volatile(68));
  FE_PHC47_map_data_volatile_28 : DEL1BWP7T port map(I => map_data_volatile(28), Z => FE_PHN47_map_data_volatile_28);
  FE_PHC46_spi_com_MISO_shift_4 : DEL1BWP7T port map(I => FE_PHN46_spi_com_MISO_shift_4, Z => spi_com_MISO_shift(4));
  FE_PHC45_map_data_volatile_59 : DEL1BWP7T port map(I => map_data_volatile(59), Z => FE_PHN45_map_data_volatile_59);
  FE_PHC44_spi_com_MISO_shift_21 : DEL1BWP7T port map(I => FE_PHN44_spi_com_MISO_shift_21, Z => spi_com_MISO_shift(21));
  FE_PHC43_map_data_volatile_19 : DEL1BWP7T port map(I => map_data_volatile(19), Z => FE_PHN43_map_data_volatile_19);
  FE_PHC42_spi_com_MISO_shift_60 : DEL1BWP7T port map(I => FE_PHN42_spi_com_MISO_shift_60, Z => spi_com_MISO_shift(60));
  FE_PHC41_map_data_volatile_27 : DEL1BWP7T port map(I => map_data_volatile(27), Z => FE_PHN41_map_data_volatile_27);
  FE_PHC40_spi_com_MISO_shift_29 : DEL1BWP7T port map(I => spi_com_MISO_shift(29), Z => FE_PHN40_spi_com_MISO_shift_29);
  FE_PHC39_map_data_volatile_64 : DEL1BWP7T port map(I => map_data_volatile(64), Z => FE_PHN39_map_data_volatile_64);
  FE_PHC38_map_data_volatile_60 : DEL1BWP7T port map(I => FE_PHN38_map_data_volatile_60, Z => map_data_volatile(60));
  FE_PHC37_spi_com_MISO_shift_54 : DEL1BWP7T port map(I => spi_com_MISO_shift(54), Z => FE_PHN37_spi_com_MISO_shift_54);
  FE_PHC36_map_data_volatile_13 : DEL1BWP7T port map(I => FE_PHN36_map_data_volatile_13, Z => map_data_volatile(13));
  FE_PHC35_spi_com_MISO_shift_22 : DEL1BWP7T port map(I => spi_com_MISO_shift(22), Z => FE_PHN35_spi_com_MISO_shift_22);
  FE_PHC34_spi_com_MISO_shift_19 : DEL1BWP7T port map(I => FE_PHN34_spi_com_MISO_shift_19, Z => spi_com_MISO_shift(19));
  FE_PHC33_map_data_volatile_65 : DEL1BWP7T port map(I => map_data_volatile(65), Z => FE_PHN33_map_data_volatile_65);
  FE_PHC32_spi_com_MISO_shift_67 : DEL1BWP7T port map(I => spi_com_MISO_shift(67), Z => FE_PHN32_spi_com_MISO_shift_67);
  FE_PHC31_spi_com_MISO_shift_48 : DEL1BWP7T port map(I => FE_PHN31_spi_com_MISO_shift_48, Z => spi_com_MISO_shift(48));
  FE_PHC30_spi_com_MISO_shift_15 : DEL1BWP7T port map(I => spi_com_MISO_shift(15), Z => FE_PHN30_spi_com_MISO_shift_15);
  FE_PHC29_spi_com_MISO_shift_31 : DEL1BWP7T port map(I => spi_com_MISO_shift(31), Z => FE_PHN29_spi_com_MISO_shift_31);
  FE_PHC28_spi_com_MISO_shift_68 : DEL1BWP7T port map(I => spi_com_MISO_shift(68), Z => FE_PHN28_spi_com_MISO_shift_68);
  FE_PHC27_spi_com_MISO_shift_23 : DEL1BWP7T port map(I => spi_com_MISO_shift(23), Z => FE_PHN27_spi_com_MISO_shift_23);
  FE_PHC26_spi_com_MISO_shift_59 : DEL1BWP7T port map(I => spi_com_MISO_shift(59), Z => FE_PHN26_spi_com_MISO_shift_59);
  FE_PHC25_spi_com_MISO_shift_38 : DEL1BWP7T port map(I => FE_PHN25_spi_com_MISO_shift_38, Z => spi_com_MISO_shift(38));
  FE_PHC24_spi_com_MISO_shift_71 : DEL1BWP7T port map(I => spi_com_MISO_shift(71), Z => FE_PHN24_spi_com_MISO_shift_71);
  FE_PHC23_spi_com_MISO_shift_24 : DEL1BWP7T port map(I => FE_PHN23_spi_com_MISO_shift_24, Z => spi_com_MISO_shift(24));
  FE_PHC22_spi_com_MISO_shift_7 : DEL1BWP7T port map(I => FE_PHN22_spi_com_MISO_shift_7, Z => spi_com_MISO_shift(7));
  FE_PHC21_spi_com_MISO_shift_70 : DEL1BWP7T port map(I => FE_PHN21_spi_com_MISO_shift_70, Z => spi_com_MISO_shift(70));
  FE_PHC20_spi_com_MISO_shift_36 : DEL1BWP7T port map(I => spi_com_MISO_shift(36), Z => FE_PHN20_spi_com_MISO_shift_36);
  FE_PHC19_spi_com_MISO_shift_30 : DEL1BWP7T port map(I => FE_PHN19_spi_com_MISO_shift_30, Z => spi_com_MISO_shift(30));
  FE_PHC18_spi_com_MISO_shift_2 : DEL1BWP7T port map(I => FE_PHN18_spi_com_MISO_shift_2, Z => spi_com_MISO_shift(2));
  FE_PHC17_vga_com_texture_module_n_20 : DEL0BWP7T port map(I => vga_com_texture_module_n_20, Z => FE_PHN17_vga_com_texture_module_n_20);
  FE_PHC16_spi_com_MISO_shift_66 : DEL1BWP7T port map(I => FE_PHN16_spi_com_MISO_shift_66, Z => spi_com_MISO_shift(66));
  FE_PHC15_spi_com_MISO_shift_53 : DEL1BWP7T port map(I => FE_PHN15_spi_com_MISO_shift_53, Z => spi_com_MISO_shift(53));
  FE_PHC14_spi_com_MISO_shift_56 : DEL1BWP7T port map(I => spi_com_MISO_shift(56), Z => FE_PHN14_spi_com_MISO_shift_56);
  FE_PHC13_spi_com_MISO_shift_69 : DEL1BWP7T port map(I => spi_com_MISO_shift(69), Z => FE_PHN13_spi_com_MISO_shift_69);
  FE_PHC12_spi_com_MISO_shift_8 : DEL1BWP7T port map(I => spi_com_MISO_shift(8), Z => FE_PHN12_spi_com_MISO_shift_8);
  FE_PHC11_spi_com_MISO_shift_37 : DEL1BWP7T port map(I => FE_PHN11_spi_com_MISO_shift_37, Z => spi_com_MISO_shift(37));
  FE_PHC10_spi_com_MISO_shift_16 : DEL1BWP7T port map(I => spi_com_MISO_shift(16), Z => FE_PHN10_spi_com_MISO_shift_16);
  FE_PHC9_spi_com_MISO_shift_63 : DEL1BWP7T port map(I => spi_com_MISO_shift(63), Z => FE_PHN9_spi_com_MISO_shift_63);
  FE_PHC8_spi_com_MISO_shift_5 : DEL1BWP7T port map(I => spi_com_MISO_shift(5), Z => FE_PHN8_spi_com_MISO_shift_5);
  FE_PDC7_vga_com_tile_module_n_914 : DEL01BWP7T port map(I => vga_com_tile_module_n_914, Z => FE_PDN7_vga_com_tile_module_n_914);
  FE_OFC6_spi_com_n_131 : DEL01BWP7T port map(I => spi_com_n_131, Z => FE_OFN6_spi_com_n_131);
  FE_OFC5_spi_com_n_139 : DEL01BWP7T port map(I => spi_com_n_139, Z => FE_OFN5_spi_com_n_139);
  FE_OFC4_vga_com_row_2 : BUFFD1P5BWP7T port map(I => vga_com_row(2), Z => FE_OFN4_vga_com_row_2);
  FE_OFC3_vga_com_row_1 : BUFFD1P5BWP7T port map(I => vga_com_row(1), Z => FE_OFN3_vga_com_row_1);
  FE_OFC2_vga_com_tile_address_0 : BUFFD1P5BWP7T port map(I => vga_com_tile_address(0), Z => FE_OFN2_vga_com_tile_address_0);
  FE_OFC1_vga_com_row_0 : BUFFD2BWP7T port map(I => vga_com_row(0), Z => FE_OFN1_vga_com_row_0);
  FE_OFC0_reset : BUFFD1P5BWP7T port map(I => reset, Z => FE_OFN0_reset);
  CTS_ccl_a_BUF_clk_G0_L2_5 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_23);
  CTS_ccl_a_BUF_clk_G0_L2_4 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_22);
  CTS_ccl_a_BUF_clk_G0_L2_3 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_21);
  CTS_ccl_a_BUF_clk_G0_L2_2 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_20);
  CTS_ccl_a_BUF_clk_G0_L2_1 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_19);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD10BWP7T port map(I => clk, Z => CTS_24);
  FE_DBTC0_reset : INVD2BWP7T port map(I => FE_OFN0_reset, ZN => FE_DBTN0_reset);
  vga_com_display_controller_module_display_state_reg_0 : DFQD0BWP7T port map(CP => CTS_23, D => n_142, Q => vga_com_display_controller_module_display_state(0));
  vga_com_display_controller_module_hsync_state_reg_0 : DFQD0BWP7T port map(CP => CTS_23, D => n_143, Q => n_116);
  g1316 : INVD5BWP7T port map(I => n_116, ZN => hsync);
  g1320 : IINR4D0BWP7T port map(A1 => FE_PHN235_vga_com_hcount_9, A2 => FE_PHN161_vga_com_hcount_7, B1 => n_106, B2 => vga_com_hcount(8), ZN => n_112);
  g1321 : MOAI22D0BWP7T port map(A1 => n_102, A2 => n_99, B1 => n_108, B2 => FE_PHN235_vga_com_hcount_9, ZN => n_111);
  vga_com_display_controller_module_vsync_state_reg_0 : DFQD1BWP7T port map(CP => CTS_23, D => n_109, Q => n_110);
  g1323 : INVD5BWP7T port map(I => n_110, ZN => vsync);
  g1324 : NR2XD0BWP7T port map(A1 => FE_PHN333_n_144, A2 => FE_OFN0_reset, ZN => n_109);
  g1325 : AO21D0BWP7T port map(A1 => n_105, A2 => vga_com_hcount(7), B => vga_com_hcount(8), Z => n_108);
  g1327 : AOI21D0BWP7T port map(A1 => n_103, A2 => vga_com_hcount(5), B => n_104, ZN => n_106);
  g1328 : OR4D1BWP7T port map(A1 => vga_com_hcount(0), A2 => vga_com_hcount(1), A3 => vga_com_hcount(2), A4 => n_100, Z => n_105);
  g1329 : MUX2ND0BWP7T port map(I0 => n_103, I1 => vga_com_hcount(5), S => vga_com_hcount(6), ZN => n_104);
  g1330 : AOI31D0BWP7T port map(A1 => n_98, A2 => vga_com_hcount(1), A3 => vga_com_hcount(0), B => vga_com_hcount(4), ZN => n_103);
  g1331 : NR4D0BWP7T port map(A1 => n_97, A2 => vga_com_vcount(3), A3 => vga_com_vcount(1), A4 => vga_com_vcount(0), ZN => n_102);
  g1332 : NR3D0BWP7T port map(A1 => n_99, A2 => n_97, A3 => FE_PHN241_vga_com_vcount_9, ZN => n_101);
  g1333 : OR4D1BWP7T port map(A1 => vga_com_hcount(3), A2 => vga_com_hcount(4), A3 => vga_com_hcount(6), A4 => vga_com_hcount(5), Z => n_100);
  g1334 : ND4D0BWP7T port map(A1 => FE_PHN239_vga_com_vcount_8, A2 => vga_com_vcount(5), A3 => vga_com_vcount(6), A4 => FE_PHN238_vga_com_vcount_7, ZN => n_99);
  g1335 : AN2D0BWP7T port map(A1 => vga_com_hcount(2), A2 => vga_com_hcount(3), Z => n_98);
  g1336 : OR2D1BWP7T port map(A1 => dir_mined(2), A2 => MOSI_data(13), Z => send);
  g1337 : OR2D1BWP7T port map(A1 => vga_com_vcount(4), A2 => FE_PHN231_vga_com_vcount_2, Z => n_97);
  g1857 : OAI31D0BWP7T port map(A1 => n_39, A2 => n_69, A3 => n_71, B => n_29, ZN => n_84);
  g1858 : OAI31D0BWP7T port map(A1 => n_25, A2 => n_68, A3 => n_72, B => n_30, ZN => n_83);
  g1859 : OAI31D0BWP7T port map(A1 => n_27, A2 => n_67, A3 => n_70, B => n_16, ZN => n_82);
  g1860 : MOAI22D0BWP7T port map(A1 => n_70, A2 => n_43, B1 => FE_PHN160_n_89, B2 => FE_OFN0_reset, ZN => n_81);
  g1861 : MOAI22D0BWP7T port map(A1 => n_71, A2 => n_41, B1 => n_85, B2 => FE_OFN0_reset, ZN => n_80);
  g1862 : MOAI22D0BWP7T port map(A1 => n_72, A2 => n_42, B1 => FE_PHN186_n_93, B2 => FE_OFN0_reset, ZN => n_79);
  g1863 : MOAI22D0BWP7T port map(A1 => n_72, A2 => n_145, B1 => n_94, B2 => FE_OFN0_reset, ZN => n_78);
  g1864 : MOAI22D0BWP7T port map(A1 => n_72, A2 => n_65, B1 => FE_PHN201_n_95, B2 => FE_OFN0_reset, ZN => n_77);
  g1865 : MOAI22D0BWP7T port map(A1 => n_71, A2 => n_56, B1 => FE_PHN169_n_86, B2 => FE_OFN0_reset, ZN => n_76);
  g1866 : MOAI22D0BWP7T port map(A1 => n_70, A2 => n_146, B1 => FE_PHN166_n_90, B2 => FE_OFN0_reset, ZN => n_75);
  g1867 : MOAI22D0BWP7T port map(A1 => n_70, A2 => n_64, B1 => FE_PHN168_n_91, B2 => FE_OFN0_reset, ZN => n_74);
  g1868 : MOAI22D0BWP7T port map(A1 => n_71, A2 => n_66, B1 => n_87, B2 => FE_OFN0_reset, ZN => n_73);
  g1869 : OAI221D0BWP7T port map(A1 => n_60, A2 => n_26, B1 => vga_com_in_red(3), B2 => n_12, C => n_34, ZN => n_72);
  g1870 : OAI221D0BWP7T port map(A1 => n_61, A2 => n_40, B1 => vga_com_in_blue(3), B2 => n_12, C => n_34, ZN => n_71);
  g1871 : OAI221D0BWP7T port map(A1 => n_62, A2 => n_28, B1 => vga_com_in_green(3), B2 => n_12, C => n_34, ZN => n_70);
  g1872 : AOI21D0BWP7T port map(A1 => n_63, A2 => n_37, B => n_23, ZN => n_69);
  g1873 : AOI21D0BWP7T port map(A1 => n_58, A2 => n_17, B => n_35, ZN => n_68);
  g1874 : AOI21D0BWP7T port map(A1 => n_59, A2 => n_21, B => n_24, ZN => n_67);
  g1875 : MAOI22D0BWP7T port map(A1 => n_63, A2 => n_47, B1 => n_63, B2 => n_47, ZN => n_66);
  g1876 : MAOI22D0BWP7T port map(A1 => n_58, A2 => n_48, B1 => n_58, B2 => n_48, ZN => n_65);
  g1877 : MAOI22D0BWP7T port map(A1 => n_59, A2 => n_44, B1 => n_59, B2 => n_44, ZN => n_64);
  g1878 : OA21D0BWP7T port map(A1 => n_51, A2 => n_24, B => n_21, Z => n_62);
  g1879 : OA21D0BWP7T port map(A1 => n_50, A2 => n_23, B => n_37, Z => n_61);
  g1880 : OA21D0BWP7T port map(A1 => n_52, A2 => n_35, B => n_17, Z => n_60);
  g1881 : OAI21D0BWP7T port map(A1 => n_19, A2 => n_31, B => n_22, ZN => n_63);
  g1883 : MAOI22D0BWP7T port map(A1 => n_46, A2 => n_31, B1 => n_46, B2 => n_31, ZN => n_56);
  g1885 : OAI21D0BWP7T port map(A1 => n_38, A2 => n_33, B => n_18, ZN => n_59);
  g1886 : OAI21D0BWP7T port map(A1 => n_36, A2 => n_32, B => n_20, ZN => n_58);
  g1889 : AOI21D0BWP7T port map(A1 => n_20, A2 => n_13, B => n_36, ZN => n_52);
  g1890 : AOI21D0BWP7T port map(A1 => n_18, A2 => n_14, B => n_38, ZN => n_51);
  g1891 : AOI21D0BWP7T port map(A1 => n_22, A2 => n_15, B => n_19, ZN => n_50);
  g1892 : IND2D1BWP7T port map(A1 => n_38, B1 => n_18, ZN => n_49);
  g1893 : IND2D1BWP7T port map(A1 => n_35, B1 => n_17, ZN => n_48);
  g1894 : IND2D1BWP7T port map(A1 => n_23, B1 => n_37, ZN => n_47);
  g1895 : INR2D1BWP7T port map(A1 => n_22, B1 => n_19, ZN => n_46);
  g1896 : IAO21D0BWP7T port map(A1 => vga_com_dim(0), A2 => n_14, B => n_33, ZN => n_43);
  g1897 : IAO21D0BWP7T port map(A1 => vga_com_dim(0), A2 => n_13, B => n_32, ZN => n_42);
  g1898 : IAO21D0BWP7T port map(A1 => vga_com_dim(0), A2 => n_15, B => n_31, ZN => n_41);
  g1899 : IND2D1BWP7T port map(A1 => n_36, B1 => n_20, ZN => n_45);
  g1900 : IND2D1BWP7T port map(A1 => n_24, B1 => n_21, ZN => n_44);
  g1901 : CKND1BWP7T port map(I => n_39, ZN => n_40);
  g1902 : ND2D1BWP7T port map(A1 => n_96, A2 => FE_OFN0_reset, ZN => n_30);
  g1903 : ND2D1BWP7T port map(A1 => n_88, A2 => FE_OFN0_reset, ZN => n_29);
  g1904 : ND2D1BWP7T port map(A1 => n_12, A2 => vga_com_in_blue(3), ZN => n_39);
  g1905 : INR2D1BWP7T port map(A1 => vga_com_dim(1), B1 => vga_com_in_green(1), ZN => n_38);
  g1906 : IND2D1BWP7T port map(A1 => vga_com_in_blue(2), B1 => vga_com_dim(2), ZN => n_37);
  g1907 : INR2D1BWP7T port map(A1 => vga_com_dim(1), B1 => vga_com_in_red(1), ZN => n_36);
  g1908 : INR2XD0BWP7T port map(A1 => vga_com_in_red(2), B1 => vga_com_dim(2), ZN => n_35);
  g1909 : NR2XD0BWP7T port map(A1 => FE_OFN0_reset, A2 => FE_PHN222_vga_com_display_controller_module_display_state_0, ZN => n_34);
  g1910 : INR2D1BWP7T port map(A1 => vga_com_dim(0), B1 => vga_com_in_green(0), ZN => n_33);
  g1911 : INR2D1BWP7T port map(A1 => vga_com_dim(0), B1 => vga_com_in_red(0), ZN => n_32);
  g1912 : INR2D1BWP7T port map(A1 => vga_com_dim(0), B1 => vga_com_in_blue(0), ZN => n_31);
  g1913 : CKND1BWP7T port map(I => n_27, ZN => n_28);
  g1914 : CKND1BWP7T port map(I => n_25, ZN => n_26);
  g1915 : ND2D1BWP7T port map(A1 => n_92, A2 => FE_OFN0_reset, ZN => n_16);
  g1916 : ND2D1BWP7T port map(A1 => n_12, A2 => vga_com_in_green(3), ZN => n_27);
  g1917 : ND2D1BWP7T port map(A1 => n_12, A2 => vga_com_in_red(3), ZN => n_25);
  g1918 : INR2XD0BWP7T port map(A1 => vga_com_in_green(2), B1 => vga_com_dim(2), ZN => n_24);
  g1919 : INR2XD0BWP7T port map(A1 => vga_com_in_blue(2), B1 => vga_com_dim(2), ZN => n_23);
  g1920 : IND2D1BWP7T port map(A1 => vga_com_dim(1), B1 => vga_com_in_blue(1), ZN => n_22);
  g1921 : IND2D1BWP7T port map(A1 => vga_com_in_green(2), B1 => vga_com_dim(2), ZN => n_21);
  g1922 : IND2D1BWP7T port map(A1 => vga_com_dim(1), B1 => vga_com_in_red(1), ZN => n_20);
  g1923 : INR2D1BWP7T port map(A1 => vga_com_dim(1), B1 => vga_com_in_blue(1), ZN => n_19);
  g1924 : IND2D1BWP7T port map(A1 => vga_com_dim(1), B1 => vga_com_in_green(1), ZN => n_18);
  g1925 : IND2D1BWP7T port map(A1 => vga_com_in_red(2), B1 => vga_com_dim(2), ZN => n_17);
  g1926 : INVD0BWP7T port map(I => vga_com_in_blue(0), ZN => n_15);
  g1927 : INVD0BWP7T port map(I => vga_com_in_green(0), ZN => n_14);
  g1928 : INVD0BWP7T port map(I => vga_com_in_red(0), ZN => n_13);
  g1929 : INVD1BWP7T port map(I => vga_com_dim(3), ZN => n_12);
  drc_bufs1930 : INVD5BWP7T port map(I => n_11, ZN => red(3));
  drc_bufs1934 : INVD5BWP7T port map(I => n_10, ZN => green(3));
  drc_bufs1938 : INVD5BWP7T port map(I => n_9, ZN => blue(3));
  drc_bufs1942 : INVD5BWP7T port map(I => n_8, ZN => blue(2));
  drc_bufs1946 : INVD5BWP7T port map(I => n_7, ZN => red(0));
  drc_bufs1950 : INVD5BWP7T port map(I => n_6, ZN => green(0));
  drc_bufs1954 : INVD5BWP7T port map(I => n_5, ZN => green(1));
  drc_bufs1958 : INVD5BWP7T port map(I => n_4, ZN => green(2));
  drc_bufs1962 : INVD5BWP7T port map(I => n_3, ZN => red(2));
  drc_bufs1966 : INVD5BWP7T port map(I => n_2, ZN => blue(0));
  drc_bufs1970 : INVD5BWP7T port map(I => n_1, ZN => red(1));
  drc_bufs1974 : INVD5BWP7T port map(I => n_0, ZN => blue(1));
  g2 : IAO21D0BWP7T port map(A1 => n_111, A2 => FE_PHN241_vga_com_vcount_9, B => FE_OFN0_reset, ZN => n_142);
  g1977 : INR2D1BWP7T port map(A1 => n_112, B1 => FE_OFN0_reset, ZN => n_143);
  g1978 : ND3D0BWP7T port map(A1 => n_101, A2 => vga_com_vcount(3), A3 => vga_com_vcount(1), ZN => n_144);
  g1979 : XNR2D1BWP7T port map(A1 => n_45, A2 => n_32, ZN => n_145);
  g1980 : XNR2D1BWP7T port map(A1 => n_49, A2 => n_33, ZN => n_146);
  vga_com_display_controller_module_red_reg_3 : DFD1BWP7T port map(CP => CTS_23, D => n_83, Q => FE_PHN165_n_96, QN => n_11);
  vga_com_display_controller_module_green_reg_3 : DFD1BWP7T port map(CP => CTS_23, D => n_82, Q => FE_PHN164_n_92, QN => n_10);
  vga_com_display_controller_module_blue_reg_3 : DFD1BWP7T port map(CP => CTS_23, D => n_84, Q => FE_PHN159_n_88, QN => n_9);
  vga_com_display_controller_module_blue_reg_2 : DFD1BWP7T port map(CP => CTS_23, D => n_73, Q => FE_PHN373_n_87, QN => n_8);
  vga_com_display_controller_module_red_reg_0 : DFD1BWP7T port map(CP => CTS_23, D => n_79, Q => n_93, QN => n_7);
  vga_com_display_controller_module_green_reg_0 : DFD1BWP7T port map(CP => CTS_23, D => n_81, Q => n_89, QN => n_6);
  vga_com_display_controller_module_green_reg_1 : DFD1BWP7T port map(CP => CTS_23, D => n_75, Q => n_90, QN => n_5);
  vga_com_display_controller_module_green_reg_2 : DFD1BWP7T port map(CP => CTS_23, D => n_74, Q => n_91, QN => n_4);
  vga_com_display_controller_module_red_reg_2 : DFD1BWP7T port map(CP => CTS_23, D => n_77, Q => n_95, QN => n_3);
  vga_com_display_controller_module_blue_reg_0 : DFD1BWP7T port map(CP => CTS_23, D => n_80, Q => FE_PHN163_n_85, QN => n_2);
  vga_com_display_controller_module_red_reg_1 : DFD1BWP7T port map(CP => CTS_23, D => n_78, Q => FE_PHN167_n_94, QN => n_1);
  vga_com_display_controller_module_blue_reg_1 : DFD1BWP7T port map(CP => CTS_23, D => n_76, Q => n_86, QN => n_0);
  fsm_com_g6646 : AO221D0BWP7T port map(A1 => fsm_com_n_529, A2 => fsm_com_n_550, B1 => fsm_com_n_530, B2 => fsm_com_n_548, C => fsm_com_n_535, Z => MOSI_data(13));
  fsm_com_g6647 : OR2D1BWP7T port map(A1 => fsm_com_n_558, A2 => dir_mined(1), Z => dir_mined(2));
  fsm_com_edge_detec3_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN100_fsm_com_edge_detec2_0, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec3(0));
  fsm_com_edge_detec3_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN123_fsm_com_edge_detec2_1, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec3(1));
  fsm_com_edge_detec3_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN93_fsm_com_edge_detec2_2, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec3(2));
  fsm_com_edge_detec3_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN212_fsm_com_edge_detec2_3, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec3(3));
  fsm_com_g6652 : AOI21D0BWP7T port map(A1 => fsm_com_n_531, A2 => fsm_com_n_532, B => fsm_com_n_516, ZN => fsm_com_n_535);
  fsm_com_g6653 : OAI31D0BWP7T port map(A1 => fsm_com_n_517, A2 => fsm_com_n_560, A3 => fsm_com_n_539, B => fsm_com_n_533, ZN => fsm_com_n_558);
  fsm_com_g6654 : ND2D1BWP7T port map(A1 => fsm_com_n_534, A2 => fsm_com_n_533, ZN => dir_mined(0));
  fsm_com_g6655 : IOA21D1BWP7T port map(A1 => fsm_com_n_528, A2 => fsm_com_n_555, B => fsm_com_n_534, ZN => dir_mined(1));
  fsm_com_edge_detec2_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN136_fsm_com_edge_detec1_2, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec2(2));
  fsm_com_edge_detec2_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN91_fsm_com_edge_detec1_0, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec2(0));
  fsm_com_edge_detec2_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN120_fsm_com_edge_detec1_1, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec2(1));
  fsm_com_edge_detec2_reg_3 : DFKCNQD1BWP7T port map(CN => fsm_com_edge_detec1(3), CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec2(3));
  fsm_com_g6660 : AO21D0BWP7T port map(A1 => fsm_com_n_564, A2 => fsm_com_n_525, B => fsm_com_n_560, Z => fsm_com_n_532);
  fsm_com_g6661 : AO21D0BWP7T port map(A1 => fsm_com_n_570, A2 => fsm_com_n_522, B => fsm_com_n_562, Z => fsm_com_n_531);
  fsm_com_g6662 : OAI211D1BWP7T port map(A1 => map_data(36), A2 => fsm_com_n_521, B => fsm_com_n_526, C => fsm_com_n_557, ZN => fsm_com_n_534);
  fsm_com_g6663 : AO21D0BWP7T port map(A1 => fsm_com_n_519, A2 => map_data(52), B => fsm_com_n_529, Z => fsm_com_n_539);
  fsm_com_g6664 : OAI211D1BWP7T port map(A1 => map_data(18), A2 => fsm_com_n_523, B => fsm_com_n_527, C => fsm_com_n_561, ZN => fsm_com_n_533);
  fsm_com_g6665 : IND2D1BWP7T port map(A1 => fsm_com_n_568, B1 => fsm_com_n_567, ZN => fsm_com_n_530);
  fsm_com_g6666 : MOAI22D0BWP7T port map(A1 => fsm_com_n_520, A2 => map_data(33), B1 => fsm_com_n_520, B2 => map_data(33), ZN => fsm_com_n_528);
  fsm_com_g6667 : ND2D1BWP7T port map(A1 => fsm_com_n_524, A2 => fsm_com_n_536, ZN => fsm_com_n_529);
  fsm_com_edge_detec1_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN209_fsm_com_edge_detec0_3, CP => CTS_19, D => FE_DBTN0_reset, Q => FE_PHN210_fsm_com_edge_detec1_3);
  fsm_com_edge_detec1_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN79_fsm_com_edge_detec0_1, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec1(1));
  fsm_com_edge_detec1_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN105_fsm_com_edge_detec0_0, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec1(0));
  fsm_com_edge_detec1_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN80_fsm_com_edge_detec0_2, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec1(2));
  fsm_com_g6672 : IND2D1BWP7T port map(A1 => fsm_com_n_569, B1 => map_data(33), ZN => fsm_com_n_567);
  fsm_com_g6673 : ND2D1BWP7T port map(A1 => fsm_com_n_523, A2 => map_data(18), ZN => fsm_com_n_527);
  fsm_com_g6674 : ND2D1BWP7T port map(A1 => fsm_com_n_521, A2 => map_data(36), ZN => fsm_com_n_526);
  fsm_com_g6675 : INR2D1BWP7T port map(A1 => fsm_com_n_538, B1 => fsm_com_n_543, ZN => game_state(0));
  fsm_com_g6676 : IND2D1BWP7T port map(A1 => fsm_com_n_572, B1 => map_data(18), ZN => fsm_com_n_570);
  fsm_com_g6677 : OR3XD1BWP7T port map(A1 => map_data(52), A2 => map_data(53), A3 => map_data(51), Z => fsm_com_n_536);
  fsm_com_g6678 : IND2D1BWP7T port map(A1 => fsm_com_n_566, B1 => map_data(36), ZN => fsm_com_n_564);
  fsm_com_g6679 : OR2D1BWP7T port map(A1 => fsm_com_n_545, A2 => fsm_com_n_544, Z => fsm_com_n_543);
  fsm_com_g6680 : AOI21D0BWP7T port map(A1 => fsm_com_n_518, A2 => fsm_com_n_556, B => fsm_com_n_517, ZN => game_state(1));
  fsm_com_g6681 : NR2D1BWP7T port map(A1 => fsm_com_n_517, A2 => fsm_com_n_556, ZN => fsm_com_n_546);
  fsm_com_g6682 : NR2XD0BWP7T port map(A1 => fsm_com_n_562, A2 => fsm_com_n_516, ZN => fsm_com_n_549);
  fsm_com_edge_detec0_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN195_button_up, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec0(2));
  fsm_com_edge_detec0_reg_3 : DFKCNQD1BWP7T port map(CN => button_down, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec0(3));
  fsm_com_g6685 : NR2XD0BWP7T port map(A1 => fsm_com_n_560, A2 => fsm_com_n_551, ZN => fsm_com_n_550);
  fsm_com_g6686 : NR2D1BWP7T port map(A1 => fsm_com_n_518, A2 => fsm_com_n_551, ZN => fsm_com_n_548);
  fsm_com_edge_detec0_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN207_button_left, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec0(0));
  fsm_com_g6688 : NR2XD0BWP7T port map(A1 => fsm_com_n_516, A2 => fsm_com_n_556, ZN => fsm_com_n_555);
  fsm_com_g6689 : OR2D1BWP7T port map(A1 => fsm_com_n_518, A2 => fsm_com_n_563, Z => fsm_com_n_538);
  fsm_com_g6690 : NR2XD0BWP7T port map(A1 => fsm_com_n_562, A2 => fsm_com_n_563, ZN => fsm_com_n_561);
  fsm_com_g6691 : NR2XD0BWP7T port map(A1 => fsm_com_n_562, A2 => fsm_com_n_517, ZN => fsm_com_n_557);
  fsm_com_edge_detec0_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN196_button_right, CP => CTS_19, D => FE_DBTN0_reset, Q => fsm_com_edge_detec0(1));
  fsm_com_g6693 : INVD0BWP7T port map(I => fsm_com_n_565, ZN => fsm_com_n_525);
  fsm_com_g6694 : INVD0BWP7T port map(I => fsm_com_n_524, ZN => fsm_com_n_537);
  fsm_com_g6695 : INVD0BWP7T port map(I => fsm_com_n_571, ZN => fsm_com_n_522);
  fsm_com_g6696 : NR2D1BWP7T port map(A1 => fsm_com_n_560, A2 => fsm_com_n_516, ZN => fsm_com_n_547);
  fsm_com_g6697 : CKXOR2D0BWP7T port map(A1 => map_data(51), A2 => map_data(53), Z => fsm_com_n_519);
  fsm_com_g6698 : NR2XD0BWP7T port map(A1 => fsm_com_n_560, A2 => fsm_com_n_517, ZN => fsm_com_n_559);
  fsm_com_g6699 : NR3D0BWP7T port map(A1 => map_data(37), A2 => map_data(38), A3 => map_data(36), ZN => fsm_com_n_565);
  fsm_com_g6700 : IND3D0BWP7T port map(A1 => map_data(52), B1 => map_data(53), B2 => map_data(51), ZN => fsm_com_n_524);
  fsm_com_g6701 : NR3D0BWP7T port map(A1 => map_data(34), A2 => map_data(35), A3 => map_data(33), ZN => fsm_com_n_568);
  fsm_com_g6702 : NR2XD0BWP7T port map(A1 => fsm_com_n_518, A2 => fsm_com_n_516, ZN => fsm_com_n_544);
  fsm_com_g6703 : OAI21D0BWP7T port map(A1 => fsm_com_n_514, A2 => map_data(20), B => fsm_com_n_572, ZN => fsm_com_n_523);
  fsm_com_g6704 : NR3D0BWP7T port map(A1 => map_data(19), A2 => map_data(20), A3 => map_data(18), ZN => fsm_com_n_571);
  fsm_com_g6705 : OAI21D0BWP7T port map(A1 => fsm_com_n_513, A2 => map_data(38), B => fsm_com_n_566, ZN => fsm_com_n_521);
  fsm_com_g6706 : OA21D0BWP7T port map(A1 => fsm_com_n_515, A2 => map_data(35), B => fsm_com_n_569, Z => fsm_com_n_520);
  fsm_com_g6707 : NR2XD0BWP7T port map(A1 => fsm_com_n_518, A2 => fsm_com_n_517, ZN => fsm_com_n_545);
  fsm_com_g6708 : ND2D1BWP7T port map(A1 => fsm_com_n_515, A2 => map_data(35), ZN => fsm_com_n_569);
  fsm_com_g6709 : ND2D1BWP7T port map(A1 => fsm_com_n_513, A2 => map_data(38), ZN => fsm_com_n_566);
  fsm_com_g6710 : ND2D1BWP7T port map(A1 => fsm_com_state(2), A2 => fsm_com_state(1), ZN => fsm_com_n_556);
  fsm_com_g6711 : IND2D1BWP7T port map(A1 => fsm_com_state(1), B1 => fsm_com_state(2), ZN => fsm_com_n_518);
  fsm_com_g6712 : IND2D1BWP7T port map(A1 => fsm_com_state(0), B1 => fsm_com_state(3), ZN => fsm_com_n_517);
  fsm_com_g6713 : CKND2D1BWP7T port map(A1 => fsm_com_state(3), A2 => fsm_com_state(0), ZN => fsm_com_n_563);
  fsm_com_g6714 : CKND2D1BWP7T port map(A1 => fsm_com_n_514, A2 => map_data(20), ZN => fsm_com_n_572);
  fsm_com_g6715 : OR2D1BWP7T port map(A1 => fsm_com_state(0), A2 => fsm_com_state(3), Z => fsm_com_n_551);
  fsm_com_g6716 : IND2D1BWP7T port map(A1 => fsm_com_state(2), B1 => fsm_com_state(1), ZN => fsm_com_n_560);
  fsm_com_g6717 : IND2D1BWP7T port map(A1 => fsm_com_state(3), B1 => fsm_com_state(0), ZN => fsm_com_n_516);
  fsm_com_g6718 : OR2D1BWP7T port map(A1 => fsm_com_state(2), A2 => fsm_com_state(1), Z => fsm_com_n_562);
  fsm_com_g6719 : INVD0BWP7T port map(I => map_data(34), ZN => fsm_com_n_515);
  fsm_com_g6720 : INVD0BWP7T port map(I => map_data(19), ZN => fsm_com_n_514);
  fsm_com_g6721 : INVD0BWP7T port map(I => map_data(37), ZN => fsm_com_n_513);
  fsm_com_energy_d_out_reg_3 : DFQD0BWP7T port map(CP => CTS_20, D => fsm_com_n_462, Q => energy_d(3));
  fsm_com_energy_d_out_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => fsm_com_n_486, Q => FE_PHN248_energy_d_4);
  fsm_com_energy_d_out_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => fsm_com_n_490, Q => energy_d(5));
  fsm_com_energy_d_out_reg_7 : DFQD1BWP7T port map(CP => CTS_20, D => fsm_com_n_475, Q => FE_PHN458_energy_d_7);
  fsm_com_energy_d_out_reg_8 : DFQD1BWP7T port map(CP => CTS_20, D => fsm_com_n_504, Q => FE_PHN245_energy_d_8);
  fsm_com_energy_d_out_reg_9 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN291_fsm_com_n_485, Q => energy_d(9));
  fsm_com_energy_d_out_reg_11 : DFQD1BWP7T port map(CP => CTS_20, D => fsm_com_n_484, Q => FE_PHN402_energy_d_11);
  fsm_com_energy_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN308_fsm_com_n_380, Q => fsm_com_energy(0));
  fsm_com_energy_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_597, Q => fsm_com_energy(3));
  fsm_com_energy_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_503, Q => fsm_com_energy(8));
  fsm_com_level_d_out_reg_0 : DFQD0BWP7T port map(CP => CTS_20, D => fsm_com_n_381, Q => FE_PHN250_level_d_0);
  fsm_com_level_d_out_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => fsm_com_n_338, Q => level_d(1));
  fsm_com_level_d_out_reg_2 : DFQD1BWP7T port map(CP => CTS_20, D => fsm_com_n_337, Q => level_d(2));
  fsm_com_level_d_out_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN321_fsm_com_n_340, Q => level_d(3));
  fsm_com_level_d_out_reg_4 : DFXQD1BWP7T port map(CP => CTS_20, DA => fsm_com_n_332, DB => fsm_com_n_323, Q => level_d(4), SA => FE_PHN477_level_d_4);
  fsm_com_level_d_out_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN320_fsm_com_n_359, Q => level_d(5));
  fsm_com_level_d_out_reg_6 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN329_fsm_com_n_363, Q => level_d(6));
  fsm_com_level_d_out_reg_7 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN299_fsm_com_n_357, Q => level_d(7));
  fsm_com_level_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN359_fsm_com_n_225, Q => level_abs(3));
  fsm_com_reached_high_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_606, Q => fsm_com_reached_high(0));
  fsm_com_reached_high_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_347, Q => fsm_com_reached_high(1));
  fsm_com_score_d_out_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN286_fsm_com_n_429, Q => score_d(1));
  fsm_com_score_d_out_reg_4 : DFQD0BWP7T port map(CP => CTS_22, D => fsm_com_n_443, Q => score_d(4));
  fsm_com_score_d_out_reg_6 : DFQD0BWP7T port map(CP => CTS_22, D => FE_PHN264_fsm_com_n_483, Q => score_d(6));
  fsm_com_score_d_out_reg_7 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN340_fsm_com_n_487, Q => score_d(7));
  fsm_com_score_d_out_reg_8 : DFXQD1BWP7T port map(CP => CTS_23, DA => fsm_com_n_435, DB => fsm_com_n_2, Q => score_d(8), SA => FE_PHN249_score_d_8);
  fsm_com_score_d_out_reg_9 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN296_fsm_com_n_464, Q => score_d(9));
  fsm_com_score_d_out_reg_10 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN282_fsm_com_n_466, Q => score_d(10));
  fsm_com_score_d_out_reg_11 : DFQD1BWP7T port map(CP => CTS_23, D => fsm_com_n_465, Q => score_d(11));
  fsm_com_score_d_out_reg_12 : DFXQD1BWP7T port map(CP => CTS_23, DA => fsm_com_n_450, DB => fsm_com_n_419, Q => score_d(12), SA => FE_PHN227_score_d_12);
  fsm_com_score_d_out_reg_13 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN337_fsm_com_n_473, Q => score_d(13));
  fsm_com_score_d_out_reg_14 : DFQD1BWP7T port map(CP => CTS_23, D => fsm_com_n_472, Q => score_d(14));
  fsm_com_score_d_out_reg_15 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN314_fsm_com_n_474, Q => score_d(15));
  fsm_com_state_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => fsm_com_n_510, Q => fsm_com_state(0));
  fsm_com_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_509, Q => fsm_com_state(1));
  fsm_com_state_reg_2 : DFQD1BWP7T port map(CP => CTS_19, D => fsm_com_n_511, Q => fsm_com_state(2));
  fsm_com_state_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_444, Q => fsm_com_state(3));
  fsm_com_x_pos_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_330, Q => xplayer(1));
  fsm_com_y_pos_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_400, Q => yplayer(3));
  fsm_com_g20841 : OR4D1BWP7T port map(A1 => FE_OFN0_reset, A2 => fsm_com_n_546, A3 => fsm_com_n_66, A4 => fsm_com_n_508, Z => fsm_com_n_511);
  fsm_com_g20844 : OR4D1BWP7T port map(A1 => FE_OFN0_reset, A2 => fsm_com_n_544, A3 => fsm_com_n_507, A4 => fsm_com_n_104, Z => fsm_com_n_510);
  fsm_com_g20845 : IIND4D0BWP7T port map(A1 => fsm_com_n_506, A2 => fsm_com_n_546, B1 => fsm_com_n_502, B2 => fsm_com_n_493, ZN => fsm_com_n_509);
  fsm_com_g20846 : IND4D0BWP7T port map(A1 => fsm_com_n_543, B1 => fsm_com_n_132, B2 => fsm_com_n_502, B3 => fsm_com_n_505, ZN => fsm_com_n_508);
  fsm_com_g20849 : ND4D0BWP7T port map(A1 => fsm_com_n_500, A2 => fsm_com_n_499, A3 => fsm_com_n_101, A4 => fsm_com_n_208, ZN => fsm_com_n_507);
  fsm_com_g20850 : OAI211D1BWP7T port map(A1 => fsm_com_n_0, A2 => fsm_com_n_538, B => fsm_com_n_495, C => fsm_com_n_245, ZN => fsm_com_n_506);
  fsm_com_g20851 : NR3D0BWP7T port map(A1 => fsm_com_n_496, A2 => fsm_com_n_421, A3 => fsm_com_n_220, ZN => fsm_com_n_505);
  fsm_com_g20852 : ND4D0BWP7T port map(A1 => fsm_com_n_488, A2 => fsm_com_n_115, A3 => fsm_com_n_83, A4 => FE_DBTN0_reset, ZN => fsm_com_n_504);
  fsm_com_g20853 : OAI211D1BWP7T port map(A1 => fsm_com_n_123, A2 => fsm_com_n_397, B => fsm_com_n_501, C => fsm_com_n_293, ZN => fsm_com_n_503);
  fsm_com_g20856 : AOI21D0BWP7T port map(A1 => fsm_com_n_413, A2 => fsm_com_n_221, B => fsm_com_n_498, ZN => fsm_com_n_501);
  fsm_com_g20857 : MAOI22D0BWP7T port map(A1 => fsm_com_n_145, A2 => button_mining, B1 => fsm_com_n_493, B2 => fsm_com_n_103, ZN => fsm_com_n_500);
  fsm_com_g20858 : AOI21D0BWP7T port map(A1 => fsm_com_n_492, A2 => FE_PHN363_fsm_com_n_103, B => fsm_com_n_85, ZN => fsm_com_n_502);
  fsm_com_g20865 : MAOI22D0BWP7T port map(A1 => fsm_com_n_37, A2 => fsm_com_n_0, B1 => fsm_com_n_480, B2 => fsm_com_n_92, ZN => fsm_com_n_499);
  fsm_com_g20866 : OAI221D0BWP7T port map(A1 => fsm_com_n_422, A2 => fsm_com_n_102, B1 => fsm_com_n_602, B2 => fsm_com_n_453, C => fsm_com_n_478, ZN => fsm_com_n_498);
  fsm_com_g20867 : ND4D0BWP7T port map(A1 => fsm_com_n_468, A2 => fsm_com_n_214, A3 => fsm_com_n_116, A4 => FE_DBTN0_reset, ZN => fsm_com_n_497);
  fsm_com_g20868 : OAI32D1BWP7T port map(A1 => fsm_com_n_105, A2 => fsm_com_n_93, A3 => fsm_com_n_480, B1 => fsm_com_n_537, B2 => fsm_com_n_35, ZN => fsm_com_n_496);
  fsm_com_g20869 : MAOI22D0BWP7T port map(A1 => fsm_com_n_595, A2 => fsm_com_n_46, B1 => fsm_com_n_117, B2 => fsm_com_n_162, ZN => fsm_com_n_495);
  fsm_com_g20881 : INVD0BWP7T port map(I => fsm_com_n_493, ZN => fsm_com_n_492);
  fsm_com_g20882 : OAI211D1BWP7T port map(A1 => fsm_com_n_183, A2 => fsm_com_n_437, B => fsm_com_n_461, C => fsm_com_n_367, ZN => fsm_com_n_491);
  fsm_com_g20883 : OAI211D1BWP7T port map(A1 => FE_PHN407_fsm_com_n_106, A2 => fsm_com_n_437, B => fsm_com_n_460, C => fsm_com_n_364, ZN => fsm_com_n_490);
  fsm_com_g20884 : OAI222D0BWP7T port map(A1 => fsm_com_n_448, A2 => fsm_com_n_19, B1 => fsm_com_n_183, B2 => fsm_com_n_456, C1 => fsm_com_n_177, C2 => fsm_com_n_458, ZN => fsm_com_n_489);
  fsm_com_g20885 : AOI21D0BWP7T port map(A1 => fsm_com_n_449, A2 => energy_d(8), B => fsm_com_n_471, ZN => fsm_com_n_488);
  fsm_com_g20886 : AO32D1BWP7T port map(A1 => fsm_com_n_454, A2 => score_d(6), A3 => score_d(5), B1 => fsm_com_n_470, B2 => score_d(7), Z => fsm_com_n_487);
  fsm_com_g20887 : AO211D0BWP7T port map(A1 => fsm_com_n_438, A2 => energy_d(4), B => fsm_com_n_463, C => fsm_com_n_366, Z => fsm_com_n_486);
  fsm_com_g20888 : OAI221D0BWP7T port map(A1 => fsm_com_n_456, A2 => FE_PHN407_fsm_com_n_106, B1 => fsm_com_n_112, B2 => fsm_com_n_458, C => fsm_com_n_467, ZN => fsm_com_n_485);
  fsm_com_g20889 : AO222D0BWP7T port map(A1 => fsm_com_n_457, A2 => fsm_com_n_253, B1 => fsm_com_n_449, B2 => FE_PHN410_energy_d_11, C1 => fsm_com_n_455, C2 => fsm_com_n_260, Z => fsm_com_n_484);
  fsm_com_g20890 : OAI31D0BWP7T port map(A1 => score_d(6), A2 => fsm_com_n_12, A3 => fsm_com_n_441, B => fsm_com_n_481, ZN => fsm_com_n_483);
  fsm_com_g20891 : IND3D1BWP7T port map(A1 => fsm_com_n_480, B1 => fsm_com_n_105, B2 => fsm_com_n_92, ZN => fsm_com_n_493);
  fsm_com_g20892 : ND4D0BWP7T port map(A1 => fsm_com_n_433, A2 => fsm_com_n_356, A3 => fsm_com_n_143, A4 => FE_DBTN0_reset, ZN => fsm_com_n_482);
  fsm_com_g20893 : ND2D1BWP7T port map(A1 => fsm_com_n_470, A2 => score_d(6), ZN => fsm_com_n_481);
  fsm_com_g20901 : OAI211D1BWP7T port map(A1 => fsm_com_n_382, A2 => fsm_com_n_430, B => fsm_com_n_446, C => fsm_com_n_364, ZN => fsm_com_n_479);
  fsm_com_g20902 : IOA21D0BWP7T port map(A1 => fsm_com_n_453, A2 => fsm_com_n_422, B => FE_PHN225_fsm_com_energy_8, ZN => fsm_com_n_478);
  fsm_com_g20903 : OAI22D0BWP7T port map(A1 => fsm_com_n_459, A2 => fsm_com_n_12, B1 => fsm_com_n_441, B2 => score_d(5), ZN => fsm_com_n_477);
  fsm_com_g20905 : AO222D0BWP7T port map(A1 => fsm_com_n_436, A2 => fsm_com_n_260, B1 => fsm_com_n_440, B2 => fsm_com_n_262, C1 => fsm_com_n_438, C2 => FE_PHN232_energy_d_7, Z => fsm_com_n_475);
  fsm_com_g20906 : AO22D0BWP7T port map(A1 => fsm_com_n_450, A2 => score_d(15), B1 => fsm_com_n_255, B2 => fsm_com_n_419, Z => fsm_com_n_474);
  fsm_com_g20907 : AO22D0BWP7T port map(A1 => fsm_com_n_450, A2 => score_d(13), B1 => fsm_com_n_96, B2 => fsm_com_n_419, Z => fsm_com_n_473);
  fsm_com_g20908 : AO22D0BWP7T port map(A1 => fsm_com_n_450, A2 => score_d(14), B1 => fsm_com_n_181, B2 => fsm_com_n_419, Z => FE_PHN313_fsm_com_n_472);
  fsm_com_g20909 : OAI22D0BWP7T port map(A1 => fsm_com_n_456, A2 => energy_d(0), B1 => fsm_com_n_458, B2 => energy_d(8), ZN => fsm_com_n_471);
  fsm_com_g20910 : ND3D0BWP7T port map(A1 => fsm_com_n_451, A2 => fsm_com_n_46, A3 => fsm_com_n_94, ZN => fsm_com_n_480);
  fsm_com_g20911 : OAI21D0BWP7T port map(A1 => fsm_com_n_425, A2 => fsm_com_n_303, B => fsm_com_n_447, ZN => fsm_com_n_469);
  fsm_com_g20912 : IINR4D0BWP7T port map(A1 => fsm_com_n_377, A2 => fsm_com_n_143, B1 => fsm_com_n_417, B2 => fsm_com_n_405, ZN => fsm_com_n_468);
  fsm_com_g20913 : ND2D1BWP7T port map(A1 => fsm_com_n_449, A2 => energy_d(9), ZN => fsm_com_n_467);
  fsm_com_g20914 : AO22D0BWP7T port map(A1 => fsm_com_n_435, A2 => score_d(10), B1 => fsm_com_n_182, B2 => fsm_com_n_2, Z => fsm_com_n_466);
  fsm_com_g20915 : OAI21D0BWP7T port map(A1 => fsm_com_n_424, A2 => score_d(5), B => fsm_com_n_459, ZN => fsm_com_n_470);
  fsm_com_g20917 : AO22D0BWP7T port map(A1 => fsm_com_n_435, A2 => score_d(11), B1 => fsm_com_n_254, B2 => fsm_com_n_2, Z => FE_PHN330_fsm_com_n_465);
  fsm_com_g20918 : AO22D0BWP7T port map(A1 => fsm_com_n_435, A2 => score_d(9), B1 => fsm_com_n_99, B2 => fsm_com_n_2, Z => fsm_com_n_464);
  fsm_com_g20919 : OAI22D0BWP7T port map(A1 => fsm_com_n_437, A2 => energy_d(0), B1 => fsm_com_n_439, B2 => energy_d(4), ZN => fsm_com_n_463);
  fsm_com_g20920 : MOAI22D0BWP7T port map(A1 => fsm_com_n_431, A2 => fsm_com_n_403, B1 => fsm_com_n_71, B2 => FE_PHN214_energy_d_3, ZN => fsm_com_n_462);
  fsm_com_g20921 : AOI22D0BWP7T port map(A1 => fsm_com_n_440, A2 => fsm_com_n_178, B1 => fsm_com_n_438, B2 => energy_d(6), ZN => fsm_com_n_461);
  fsm_com_g20922 : AOI22D0BWP7T port map(A1 => fsm_com_n_440, A2 => fsm_com_n_113, B1 => fsm_com_n_438, B2 => energy_d(5), ZN => fsm_com_n_460);
  fsm_com_g20923 : INVD0BWP7T port map(I => fsm_com_n_458, ZN => fsm_com_n_457);
  fsm_com_g20924 : INVD0BWP7T port map(I => fsm_com_n_455, ZN => fsm_com_n_456);
  fsm_com_g20925 : NR2XD0BWP7T port map(A1 => fsm_com_n_441, A2 => score_d(7), ZN => fsm_com_n_454);
  fsm_com_g20926 : NR2XD0BWP7T port map(A1 => fsm_com_n_442, A2 => fsm_com_n_426, ZN => fsm_com_n_459);
  fsm_com_g20927 : ND2D1BWP7T port map(A1 => fsm_com_n_436, A2 => fsm_com_n_297, ZN => fsm_com_n_458);
  fsm_com_g20928 : NR2D0BWP7T port map(A1 => fsm_com_n_437, A2 => fsm_com_n_297, ZN => fsm_com_n_455);
  fsm_com_g20934 : INVD1BWP7T port map(I => fsm_com_n_448, ZN => fsm_com_n_449);
  fsm_com_g20935 : AOI22D0BWP7T port map(A1 => fsm_com_n_420, A2 => fsm_com_n_303, B1 => fsm_com_n_71, B2 => FE_PHN403_energy_d_1, ZN => fsm_com_n_447);
  fsm_com_g20936 : AOI22D0BWP7T port map(A1 => fsm_com_n_420, A2 => fsm_com_n_382, B1 => fsm_com_n_71, B2 => FE_PHN189_energy_d_2, ZN => fsm_com_n_446);
  fsm_com_g20937 : AOI221D0BWP7T port map(A1 => fsm_com_n_261, A2 => FE_PHN206_fsm_com_energy_7, B1 => fsm_com_n_365, B2 => fsm_com_n_138, C => fsm_com_n_432, ZN => fsm_com_n_445);
  fsm_com_g20938 : OR4D1BWP7T port map(A1 => fsm_com_n_222, A2 => fsm_com_n_543, A3 => fsm_com_n_104, A4 => fsm_com_n_421, Z => fsm_com_n_444);
  fsm_com_g20939 : AO21D0BWP7T port map(A1 => fsm_com_n_426, A2 => FE_PHN244_score_d_4, B => fsm_com_n_442, Z => fsm_com_n_443);
  fsm_com_g20940 : AOI21D0BWP7T port map(A1 => fsm_com_n_210, A2 => fsm_com_n_413, B => fsm_com_n_239, ZN => fsm_com_n_453);
  fsm_com_g20941 : AOI21D0BWP7T port map(A1 => fsm_com_n_407, A2 => button_mining, B => fsm_com_n_394, ZN => fsm_com_n_451);
  fsm_com_g20942 : OR2D1BWP7T port map(A1 => fsm_com_n_435, A2 => fsm_com_n_2, Z => fsm_com_n_450);
  fsm_com_g20943 : NR2XD0BWP7T port map(A1 => fsm_com_n_440, A2 => fsm_com_n_438, ZN => fsm_com_n_448);
  fsm_com_g20944 : INVD1BWP7T port map(I => fsm_com_n_439, ZN => fsm_com_n_440);
  fsm_com_g20945 : INVD0BWP7T port map(I => fsm_com_n_437, ZN => fsm_com_n_436);
  fsm_com_g20946 : NR2XD0BWP7T port map(A1 => fsm_com_n_424, A2 => FE_PHN244_score_d_4, ZN => fsm_com_n_442);
  fsm_com_g20947 : IND2D1BWP7T port map(A1 => fsm_com_n_424, B1 => FE_PHN244_score_d_4, ZN => fsm_com_n_441);
  fsm_com_g20948 : ND2D1BWP7T port map(A1 => fsm_com_n_420, A2 => fsm_com_n_283, ZN => fsm_com_n_439);
  fsm_com_g20949 : IND2D1BWP7T port map(A1 => fsm_com_n_71, B1 => fsm_com_n_425, ZN => fsm_com_n_438);
  fsm_com_g20951 : IND2D1BWP7T port map(A1 => fsm_com_n_283, B1 => fsm_com_n_420, ZN => fsm_com_n_437);
  fsm_com_g20954 : OAI22D0BWP7T port map(A1 => fsm_com_n_3, A2 => fsm_com_n_398, B1 => fsm_com_n_115, B2 => fsm_com_n_17, ZN => fsm_com_n_434);
  fsm_com_g20955 : AOI21D0BWP7T port map(A1 => fsm_com_n_385, A2 => fsm_com_n_81, B => fsm_com_n_418, ZN => fsm_com_n_433);
  fsm_com_g20956 : AO211D0BWP7T port map(A1 => fsm_com_n_365, A2 => fsm_com_n_68, B => fsm_com_n_412, C => fsm_com_n_411, Z => fsm_com_n_432);
  fsm_com_g20957 : OA31D1BWP7T port map(A1 => fsm_com_n_151, A2 => fsm_com_n_303, A3 => fsm_com_n_382, B => fsm_com_n_425, Z => fsm_com_n_431);
  fsm_com_g20958 : OA21D0BWP7T port map(A1 => fsm_com_n_304, A2 => fsm_com_n_151, B => fsm_com_n_425, Z => fsm_com_n_430);
  fsm_com_g20959 : MOAI22D0BWP7T port map(A1 => fsm_com_n_3, A2 => fsm_com_n_307, B1 => fsm_com_n_114, B2 => FE_PHN174_score_d_1, ZN => fsm_com_n_429);
  fsm_com_g20960 : OAI22D0BWP7T port map(A1 => fsm_com_n_3, A2 => fsm_com_n_227, B1 => fsm_com_n_115, B2 => FE_PHN188_fsm_com_n_28, ZN => fsm_com_n_428);
  fsm_com_g20961 : OAI22D0BWP7T port map(A1 => fsm_com_n_3, A2 => fsm_com_n_358, B1 => fsm_com_n_115, B2 => FE_PHN184_fsm_com_n_27, ZN => fsm_com_n_427);
  fsm_com_g20962 : IND2D1BWP7T port map(A1 => fsm_com_n_426, B1 => fsm_com_n_424, ZN => fsm_com_n_435);
  fsm_com_g20963 : ND2D1BWP7T port map(A1 => fsm_com_n_596, A2 => FE_DBTN0_reset, ZN => fsm_com_n_423);
  fsm_com_g20964 : ND2D1BWP7T port map(A1 => fsm_com_n_3, A2 => fsm_com_n_115, ZN => fsm_com_n_426);
  fsm_com_g20965 : ND2D1BWP7T port map(A1 => fsm_com_n_416, A2 => fsm_com_n_152, ZN => fsm_com_n_425);
  fsm_com_g20966 : IND2D1BWP7T port map(A1 => fsm_com_n_415, B1 => fsm_com_n_166, ZN => fsm_com_n_424);
  fsm_com_g20969 : OAI211D1BWP7T port map(A1 => fsm_com_n_195, A2 => fsm_com_n_345, B => fsm_com_n_598, C => fsm_com_n_360, ZN => fsm_com_n_418);
  fsm_com_g20970 : OAI21D0BWP7T port map(A1 => fsm_com_n_383, A2 => fsm_com_n_195, B => fsm_com_n_408, ZN => fsm_com_n_417);
  fsm_com_g20971 : AO21D0BWP7T port map(A1 => fsm_com_n_397, A2 => fsm_com_n_95, B => fsm_com_n_54, Z => fsm_com_n_422);
  fsm_com_g20972 : IOA21D1BWP7T port map(A1 => fsm_com_n_394, A2 => fsm_com_n_46, B => fsm_com_n_538, ZN => fsm_com_n_421);
  fsm_com_g20973 : NR2XD0BWP7T port map(A1 => fsm_com_n_416, A2 => fsm_com_n_151, ZN => fsm_com_n_420);
  fsm_com_g20974 : NR4D0BWP7T port map(A1 => fsm_com_n_415, A2 => fsm_com_n_275, A3 => fsm_com_n_284, A4 => fsm_com_n_166, ZN => fsm_com_n_419);
  fsm_com_g20977 : AO21D0BWP7T port map(A1 => fsm_com_n_382, A2 => fsm_com_n_329, B => fsm_com_n_403, Z => fsm_com_n_416);
  fsm_com_g20978 : ND2D1BWP7T port map(A1 => fsm_com_n_402, A2 => fsm_com_n_152, ZN => fsm_com_n_415);
  fsm_com_g20982 : AOI22D0BWP7T port map(A1 => fsm_com_n_212, A2 => fsm_com_n_390, B1 => fsm_com_n_237, B2 => fsm_com_n_602, ZN => fsm_com_n_412);
  fsm_com_g20983 : OAI22D0BWP7T port map(A1 => fsm_com_n_292, A2 => fsm_com_n_390, B1 => fsm_com_n_75, B2 => fsm_com_n_23, ZN => fsm_com_n_411);
  fsm_com_g20985 : IND4D0BWP7T port map(A1 => fsm_com_n_372, B1 => fsm_com_n_290, B2 => fsm_com_n_376, B3 => fsm_com_n_388, ZN => fsm_com_n_409);
  fsm_com_g20986 : AOI211XD0BWP7T port map(A1 => fsm_com_n_139, A2 => fsm_com_energy(5), B => fsm_com_n_395, C => fsm_com_n_370, ZN => fsm_com_n_408);
  fsm_com_g20987 : IOA21D1BWP7T port map(A1 => fsm_com_n_384, A2 => FE_PHN399_fsm_com_energy_8, B => fsm_com_n_407, ZN => fsm_com_n_413);
  fsm_com_g20988 : IND3D1BWP7T port map(A1 => fsm_com_n_387, B1 => fsm_com_n_118, B2 => fsm_com_n_324, ZN => fsm_com_n_406);
  fsm_com_g20989 : AOI221D0BWP7T port map(A1 => fsm_com_n_206, A2 => fsm_com_n_383, B1 => fsm_com_n_207, B2 => fsm_com_n_26, C => fsm_com_n_80, ZN => fsm_com_n_405);
  fsm_com_g20990 : ND4D0BWP7T port map(A1 => fsm_com_n_379, A2 => fsm_com_n_137, A3 => fsm_com_n_176, A4 => FE_DBTN0_reset, ZN => fsm_com_n_404);
  fsm_com_g20991 : OR2D1BWP7T port map(A1 => fsm_com_n_384, A2 => FE_PHN456_fsm_com_energy_8, Z => fsm_com_n_407);
  fsm_com_g20994 : OAI222D0BWP7T port map(A1 => fsm_com_n_392, A2 => fsm_com_n_272, B1 => fsm_com_n_251, B2 => fsm_com_n_44, C1 => FE_PHN208_fsm_com_n_20, C2 => fsm_com_n_41, ZN => fsm_com_n_400);
  fsm_com_g20995 : MAOI22D0BWP7T port map(A1 => fsm_com_n_373, A2 => energy_d(3), B1 => fsm_com_n_373, B2 => energy_d(3), ZN => fsm_com_n_403);
  fsm_com_g20996 : AOI21D0BWP7T port map(A1 => fsm_com_n_389, A2 => fsm_com_n_307, B => fsm_com_n_398, ZN => fsm_com_n_402);
  fsm_com_g21000 : OAI222D0BWP7T port map(A1 => fsm_com_n_374, A2 => fsm_com_n_272, B1 => fsm_com_n_179, B2 => fsm_com_n_44, C1 => FE_PHN215_fsm_com_n_6, C2 => fsm_com_n_41, ZN => fsm_com_n_396);
  fsm_com_g21001 : AOI22D0BWP7T port map(A1 => fsm_com_n_212, A2 => fsm_com_n_383, B1 => fsm_com_n_238, B2 => fsm_com_n_602, ZN => fsm_com_n_395);
  fsm_com_g21002 : MOAI22D0BWP7T port map(A1 => fsm_com_n_354, A2 => fsm_com_n_17, B1 => fsm_com_n_354, B2 => fsm_com_n_17, ZN => fsm_com_n_398);
  fsm_com_g21003 : AOI21D0BWP7T port map(A1 => fsm_com_n_352, A2 => FE_PHN225_fsm_com_energy_8, B => fsm_com_n_394, ZN => fsm_com_n_397);
  fsm_com_g21004 : IND4D0BWP7T port map(A1 => fsm_com_n_346, B1 => FE_DBTN0_reset, B2 => fsm_com_n_131, B3 => fsm_com_n_137, ZN => fsm_com_n_393);
  fsm_com_g21005 : OAI222D0BWP7T port map(A1 => fsm_com_n_343, A2 => yplayer(3), B1 => yplayer(1), B2 => fsm_com_n_328, C1 => xplayer(3), C2 => fsm_com_n_270, ZN => fsm_com_n_392);
  fsm_com_g21006 : AOI22D0BWP7T port map(A1 => fsm_com_n_212, A2 => fsm_com_n_345, B1 => fsm_com_n_236, B2 => fsm_com_n_602, ZN => fsm_com_n_391);
  fsm_com_g21007 : NR2D1BWP7T port map(A1 => fsm_com_n_352, A2 => FE_PHN225_fsm_com_energy_8, ZN => fsm_com_n_394);
  fsm_com_g21010 : OAI21D0BWP7T port map(A1 => fsm_com_n_305, A2 => score_d(2), B => score_d(3), ZN => fsm_com_n_389);
  fsm_com_g21011 : OAI22D0BWP7T port map(A1 => fsm_com_n_239, A2 => fsm_com_n_368, B1 => fsm_com_n_228, B2 => FE_PHN202_fsm_com_energy_4, ZN => fsm_com_n_388);
  fsm_com_g21012 : OAI211D1BWP7T port map(A1 => fsm_com_n_58, A2 => fsm_com_n_187, B => fsm_com_n_361, C => fsm_com_n_341, ZN => fsm_com_n_387);
  fsm_com_g21013 : AOI211XD0BWP7T port map(A1 => fsm_com_n_350, A2 => FE_PHN395_fsm_com_energy_3, B => fsm_com_n_371, C => fsm_com_n_322, ZN => fsm_com_n_386);
  fsm_com_g21014 : AOI22D0BWP7T port map(A1 => fsm_com_n_345, A2 => fsm_com_n_206, B1 => fsm_com_n_207, B2 => fsm_com_n_9, ZN => fsm_com_n_385);
  fsm_com_g21015 : OA21D0BWP7T port map(A1 => fsm_com_n_333, A2 => fsm_com_n_23, B => fsm_com_n_384, Z => fsm_com_n_390);
  fsm_com_g21016 : ND2D1BWP7T port map(A1 => fsm_com_n_333, A2 => fsm_com_n_23, ZN => fsm_com_n_384);
  fsm_com_g21025 : AO211D0BWP7T port map(A1 => fsm_com_n_152, A2 => level_d(0), B => fsm_com_n_339, C => fsm_com_n_71, Z => fsm_com_n_381);
  fsm_com_g21026 : IND4D0BWP7T port map(A1 => fsm_com_n_322, B1 => fsm_com_n_116, B2 => fsm_com_n_321, B3 => fsm_com_n_308, ZN => fsm_com_n_380);
  fsm_com_g21027 : OAI211D1BWP7T port map(A1 => xplayer(1), A2 => fsm_com_n_270, B => fsm_com_n_344, C => fsm_com_n_271, ZN => fsm_com_n_379);
  fsm_com_g21028 : OAI211D1BWP7T port map(A1 => fsm_com_n_151, A2 => fsm_com_n_231, B => fsm_com_n_364, C => fsm_com_n_111, ZN => FE_PHN336_fsm_com_n_378);
  fsm_com_g21029 : AOI22D0BWP7T port map(A1 => fsm_com_n_336, A2 => fsm_com_n_68, B1 => fsm_com_n_204, B2 => fsm_com_energy(5), ZN => fsm_com_n_377);
  fsm_com_g21030 : AOI21D0BWP7T port map(A1 => fsm_com_n_273, A2 => fsm_com_n_205, B => fsm_com_n_362, ZN => fsm_com_n_376);
  fsm_com_g21031 : AOI211XD0BWP7T port map(A1 => fsm_com_n_550, A2 => fsm_com_n_557, B => fsm_com_n_349, C => fsm_com_n_327, ZN => fsm_com_n_375);
  fsm_com_g21032 : OAI222D0BWP7T port map(A1 => fsm_com_n_325, A2 => yplayer(2), B1 => yplayer(1), B2 => fsm_com_n_311, C1 => xplayer(2), C2 => fsm_com_n_270, ZN => fsm_com_n_374);
  fsm_com_g21033 : OA21D0BWP7T port map(A1 => fsm_com_n_351, A2 => fsm_com_n_26, B => fsm_com_n_314, Z => fsm_com_n_383);
  fsm_com_g21034 : OA21D0BWP7T port map(A1 => fsm_com_n_599, A2 => fsm_com_n_13, B => fsm_com_n_373, Z => fsm_com_n_382);
  fsm_com_g21035 : OAI221D0BWP7T port map(A1 => fsm_com_n_158, A2 => fsm_com_n_289, B1 => fsm_com_reached_high(1), B2 => fsm_com_n_116, C => fsm_com_n_277, ZN => fsm_com_n_372);
  fsm_com_g21036 : OAI211D1BWP7T port map(A1 => fsm_com_n_240, A2 => fsm_com_n_67, B => fsm_com_n_316, C => fsm_com_n_288, ZN => fsm_com_n_371);
  fsm_com_g21037 : AOI22D0BWP7T port map(A1 => fsm_com_n_334, A2 => fsm_com_n_268, B1 => fsm_com_n_73, B2 => fsm_com_n_119, ZN => fsm_com_n_370);
  fsm_com_g21038 : ND3D0BWP7T port map(A1 => fsm_com_n_317, A2 => fsm_com_n_137, A3 => FE_DBTN0_reset, ZN => fsm_com_n_369);
  fsm_com_g21039 : NR2D0BWP7T port map(A1 => fsm_com_n_209, A2 => fsm_com_n_355, ZN => fsm_com_n_368);
  fsm_com_g21040 : ND2D1BWP7T port map(A1 => fsm_com_n_599, A2 => fsm_com_n_13, ZN => fsm_com_n_373);
  fsm_com_g21046 : INVD0BWP7T port map(I => fsm_com_n_366, ZN => fsm_com_n_367);
  fsm_com_g21047 : AO22D0BWP7T port map(A1 => fsm_com_n_323, A2 => fsm_com_n_184, B1 => level_d(6), B2 => fsm_com_n_332, Z => fsm_com_n_363);
  fsm_com_g21048 : IAO21D0BWP7T port map(A1 => fsm_com_n_273, A2 => fsm_com_n_189, B => fsm_com_n_355, ZN => fsm_com_n_362);
  fsm_com_g21049 : AOI221D0BWP7T port map(A1 => fsm_com_n_300, A2 => fsm_com_n_91, B1 => fsm_com_n_249, B2 => fsm_com_n_242, C => fsm_com_n_600, ZN => fsm_com_n_361);
  fsm_com_g21050 : MAOI22D0BWP7T port map(A1 => fsm_com_n_204, A2 => fsm_com_energy(6), B1 => fsm_com_n_315, B2 => fsm_com_n_67, ZN => fsm_com_n_360);
  fsm_com_g21051 : AO22D0BWP7T port map(A1 => fsm_com_n_323, A2 => fsm_com_n_98, B1 => level_d(5), B2 => fsm_com_n_332, Z => fsm_com_n_359);
  fsm_com_g21052 : MAOI22D0BWP7T port map(A1 => fsm_com_n_305, A2 => FE_PHN184_fsm_com_n_27, B1 => fsm_com_n_305, B2 => FE_PHN184_fsm_com_n_27, ZN => fsm_com_n_358);
  fsm_com_g21053 : AO22D0BWP7T port map(A1 => fsm_com_n_323, A2 => fsm_com_n_256, B1 => level_d(7), B2 => fsm_com_n_332, Z => fsm_com_n_357);
  fsm_com_g21054 : AOI22D0BWP7T port map(A1 => fsm_com_n_138, A2 => fsm_com_n_335, B1 => fsm_com_n_139, B2 => fsm_com_energy(6), ZN => fsm_com_n_356);
  fsm_com_g21055 : MOAI22D0BWP7T port map(A1 => fsm_com_n_324, A2 => FE_OFN0_reset, B1 => fsm_com_n_114, B2 => FE_PHN205_fsm_com_reached_high_1, ZN => fsm_com_n_366);
  fsm_com_g21056 : OAI21D0BWP7T port map(A1 => fsm_com_n_295, A2 => fsm_com_n_23, B => fsm_com_n_352, ZN => fsm_com_n_365);
  fsm_com_g21057 : AOI22D0BWP7T port map(A1 => fsm_com_n_322, A2 => FE_DBTN0_reset, B1 => fsm_com_n_114, B2 => FE_PHN224_fsm_com_reached_high_0, ZN => fsm_com_n_364);
  fsm_com_g21058 : HA1D0BWP7T port map(A => fsm_com_n_24, B => fsm_com_n_243, CO => fsm_com_n_351, S => fsm_com_n_355);
  fsm_com_g21059 : AO221D0BWP7T port map(A1 => fsm_com_n_69, A2 => fsm_com_n_252, B1 => fsm_com_n_138, B2 => fsm_com_n_164, C => fsm_com_n_261, Z => fsm_com_n_350);
  fsm_com_g21060 : OAI211D1BWP7T port map(A1 => fsm_com_n_102, A2 => fsm_com_n_258, B => fsm_com_n_326, C => fsm_com_n_601, ZN => fsm_com_n_349);
  fsm_com_g21062 : ND2D1BWP7T port map(A1 => fsm_com_n_318, A2 => fsm_com_n_324, ZN => fsm_com_n_347);
  fsm_com_g21063 : OAI22D0BWP7T port map(A1 => fsm_com_n_306, A2 => fsm_com_n_64, B1 => fsm_com_n_230, B2 => fsm_com_n_40, ZN => fsm_com_n_346);
  fsm_com_g21064 : ND2D1BWP7T port map(A1 => fsm_com_n_305, A2 => score_d(2), ZN => fsm_com_n_354);
  fsm_com_g21066 : ND2D1BWP7T port map(A1 => fsm_com_n_295, A2 => fsm_com_n_23, ZN => fsm_com_n_352);
  fsm_com_g21068 : OAI22D0BWP7T port map(A1 => fsm_com_n_306, A2 => yplayer(1), B1 => fsm_com_n_294, B2 => FE_PHN223_fsm_com_n_8, ZN => fsm_com_n_344);
  fsm_com_g21069 : OA21D0BWP7T port map(A1 => fsm_com_n_266, A2 => fsm_com_n_10, B => fsm_com_n_325, Z => fsm_com_n_343);
  fsm_com_g21070 : OAI22D0BWP7T port map(A1 => fsm_com_n_312, A2 => FE_PHN208_fsm_com_n_20, B1 => fsm_com_n_278, B2 => xplayer(3), ZN => fsm_com_n_342);
  fsm_com_g21071 : AOI221D0BWP7T port map(A1 => fsm_com_n_72, A2 => fsm_com_n_144, B1 => fsm_com_n_55, B2 => fsm_com_energy(1), C => fsm_com_n_302, ZN => fsm_com_n_341);
  fsm_com_g21072 : MOAI22D0BWP7T port map(A1 => fsm_com_n_313, A2 => fsm_com_n_259, B1 => fsm_com_n_152, B2 => level_d(3), ZN => fsm_com_n_340);
  fsm_com_g21073 : MOAI22D0BWP7T port map(A1 => fsm_com_n_313, A2 => level_d(0), B1 => fsm_com_n_544, B2 => FE_DBTN0_reset, ZN => fsm_com_n_339);
  fsm_com_g21074 : MOAI22D0BWP7T port map(A1 => fsm_com_n_313, A2 => fsm_com_n_100, B1 => fsm_com_n_152, B2 => FE_PHN498_level_d_1, ZN => fsm_com_n_338);
  fsm_com_g21075 : MOAI22D0BWP7T port map(A1 => fsm_com_n_313, A2 => fsm_com_n_185, B1 => fsm_com_n_152, B2 => level_d(2), ZN => FE_PHN266_fsm_com_n_337);
  fsm_com_g21076 : ND2D1BWP7T port map(A1 => fsm_com_n_334, A2 => fsm_com_n_268, ZN => fsm_com_n_336);
  fsm_com_g21077 : AOI21D0BWP7T port map(A1 => fsm_com_n_314, A2 => fsm_com_energy(6), B => fsm_com_n_333, ZN => fsm_com_n_345);
  fsm_com_g21078 : INVD0BWP7T port map(I => fsm_com_n_315, ZN => fsm_com_n_335);
  fsm_com_g21079 : AO211D0BWP7T port map(A1 => fsm_com_n_269, A2 => xplayer(0), B => fsm_com_n_247, C => fsm_com_n_130, Z => fsm_com_n_331);
  fsm_com_g21080 : ND2D1BWP7T port map(A1 => fsm_com_n_274, A2 => fsm_com_energy(5), ZN => fsm_com_n_334);
  fsm_com_g21081 : AO21D0BWP7T port map(A1 => fsm_com_n_276, A2 => xplayer(1), B => fsm_com_n_301, Z => fsm_com_n_330);
  fsm_com_g21082 : IND2D1BWP7T port map(A1 => fsm_com_n_231, B1 => fsm_com_n_304, ZN => fsm_com_n_329);
  fsm_com_g21083 : ND3D0BWP7T port map(A1 => fsm_com_n_294, A2 => fsm_com_n_10, A3 => yplayer(3), ZN => fsm_com_n_328);
  fsm_com_g21084 : OA31D1BWP7T port map(A1 => fsm_com_n_42, A2 => fsm_com_n_219, A3 => fsm_com_n_250, B => FE_PHN230_fsm_com_energy_2, Z => fsm_com_n_327);
  fsm_com_g21085 : OAI31D0BWP7T port map(A1 => fsm_com_n_257, A2 => fsm_com_n_239, A3 => fsm_com_n_248, B => fsm_com_energy(2), ZN => fsm_com_n_326);
  fsm_com_g21086 : NR2D1BWP7T port map(A1 => fsm_com_n_314, A2 => fsm_com_energy(6), ZN => fsm_com_n_333);
  fsm_com_g21087 : ND2D1BWP7T port map(A1 => fsm_com_n_151, A2 => fsm_com_n_313, ZN => fsm_com_n_332);
  fsm_com_g21088 : AO31D1BWP7T port map(A1 => fsm_com_n_602, A2 => fsm_com_n_264, A3 => fsm_com_n_158, B => fsm_com_energy(0), Z => fsm_com_n_321);
  fsm_com_g21089 : AOI22D0BWP7T port map(A1 => fsm_com_n_265, A2 => fsm_com_n_252, B1 => fsm_com_n_138, B2 => fsm_com_n_241, ZN => fsm_com_n_320);
  fsm_com_g21091 : OAI21D0BWP7T port map(A1 => fsm_com_n_286, A2 => fsm_com_n_545, B => FE_PHN205_fsm_com_reached_high_1, ZN => fsm_com_n_318);
  fsm_com_g21092 : OA22D0BWP7T port map(A1 => fsm_com_n_296, A2 => FE_PHN215_fsm_com_n_6, B1 => xplayer(2), B2 => fsm_com_n_291, Z => fsm_com_n_317);
  fsm_com_g21093 : OAI22D0BWP7T port map(A1 => fsm_com_n_235, A2 => fsm_com_n_228, B1 => fsm_com_n_211, B2 => fsm_com_n_252, ZN => fsm_com_n_316);
  fsm_com_g21094 : IAO21D0BWP7T port map(A1 => fsm_com_n_266, A2 => fsm_com_n_8, B => fsm_com_n_306, ZN => fsm_com_n_325);
  fsm_com_g21095 : OAI21D0BWP7T port map(A1 => fsm_com_n_282, A2 => fsm_com_n_192, B => fsm_com_n_545, ZN => fsm_com_n_324);
  fsm_com_g21096 : AOI211XD0BWP7T port map(A1 => fsm_com_n_226, A2 => fsm_com_n_256, B => fsm_com_n_285, C => fsm_com_n_115, ZN => fsm_com_n_323);
  fsm_com_g21097 : OA21D0BWP7T port map(A1 => fsm_com_n_232, A2 => fsm_com_n_282, B => fsm_com_n_545, Z => fsm_com_n_322);
  fsm_com_g21098 : OA221D0BWP7T port map(A1 => fsm_com_n_29, A2 => xplayer(2), B1 => FE_PHN215_fsm_com_n_6, B2 => fsm_com_n_35, C => fsm_com_n_296, Z => fsm_com_n_312);
  fsm_com_g21099 : ND2D0BWP7T port map(A1 => fsm_com_n_294, A2 => yplayer(2), ZN => fsm_com_n_311);
  fsm_com_g21100 : NR2D1BWP7T port map(A1 => fsm_com_n_214, A2 => fsm_com_n_282, ZN => fsm_com_n_310);
  fsm_com_g21101 : AOI21D0BWP7T port map(A1 => fsm_com_n_215, A2 => fsm_com_n_7, B => dir_mined(2), ZN => fsm_com_n_309);
  fsm_com_g21102 : OAI31D0BWP7T port map(A1 => fsm_com_n_242, A2 => fsm_com_n_246, A3 => fsm_com_n_239, B => FE_PHN397_fsm_com_energy_0, ZN => fsm_com_n_308);
  fsm_com_g21103 : AOI21D0BWP7T port map(A1 => fsm_com_n_268, A2 => fsm_com_energy(6), B => fsm_com_n_295, ZN => fsm_com_n_315);
  fsm_com_g21104 : ND2D1BWP7T port map(A1 => fsm_com_n_243, A2 => fsm_com_n_84, ZN => fsm_com_n_314);
  fsm_com_g21105 : ND2D1BWP7T port map(A1 => fsm_com_n_285, A2 => fsm_com_n_114, ZN => fsm_com_n_313);
  fsm_com_g21106 : INVD0BWP7T port map(I => fsm_com_n_304, ZN => fsm_com_n_303);
  fsm_com_g21107 : AOI211D1BWP7T port map(A1 => fsm_com_n_224, A2 => fsm_com_n_91, B => fsm_com_n_198, C => fsm_com_n_200, ZN => fsm_com_n_302);
  fsm_com_g21108 : OAI31D0BWP7T port map(A1 => xplayer(1), A2 => FE_PHN233_fsm_com_n_22, A3 => fsm_com_n_73, B => fsm_com_n_281, ZN => fsm_com_n_301);
  fsm_com_g21109 : AO211D0BWP7T port map(A1 => fsm_com_n_249, A2 => fsm_com_n_69, B => fsm_com_n_244, C => fsm_com_n_228, Z => fsm_com_n_300);
  fsm_com_g21110 : MAOI22D0BWP7T port map(A1 => fsm_com_n_265, A2 => fsm_com_n_180, B1 => fsm_com_n_123, B2 => fsm_com_n_186, ZN => fsm_com_n_299);
  fsm_com_g21111 : MOAI22D0BWP7T port map(A1 => fsm_com_n_223, A2 => fsm_com_n_65, B1 => fsm_com_n_137, B2 => level_abs(4), ZN => fsm_com_n_298);
  fsm_com_g21112 : MAOI22D0BWP7T port map(A1 => fsm_com_n_233, A2 => fsm_com_n_216, B1 => fsm_com_n_233, B2 => fsm_com_n_216, ZN => fsm_com_n_307);
  fsm_com_g21113 : OAI21D0BWP7T port map(A1 => fsm_com_n_266, A2 => fsm_com_n_11, B => fsm_com_n_548, ZN => fsm_com_n_306);
  fsm_com_g21114 : OAI21D0BWP7T port map(A1 => fsm_com_n_218, A2 => fsm_com_n_216, B => fsm_com_n_217, ZN => fsm_com_n_305);
  fsm_com_g21115 : MOAI22D0BWP7T port map(A1 => fsm_com_n_97, A2 => fsm_com_n_215, B1 => fsm_com_n_97, B2 => fsm_com_n_215, ZN => fsm_com_n_304);
  fsm_com_g21116 : OAI31D0BWP7T port map(A1 => fsm_com_n_42, A2 => fsm_com_n_204, A3 => fsm_com_n_199, B => FE_PHN225_fsm_com_energy_8, ZN => fsm_com_n_293);
  fsm_com_g21117 : AOI21D0BWP7T port map(A1 => fsm_com_n_69, A2 => fsm_com_energy(7), B => fsm_com_n_265, ZN => fsm_com_n_292);
  fsm_com_g21118 : AOI21D0BWP7T port map(A1 => fsm_com_n_234, A2 => fsm_com_n_550, B => fsm_com_n_122, ZN => fsm_com_n_291);
  fsm_com_g21119 : OAI21D0BWP7T port map(A1 => fsm_com_n_232, A2 => fsm_com_n_192, B => fsm_com_n_545, ZN => fsm_com_n_290);
  fsm_com_g21120 : OA21D0BWP7T port map(A1 => fsm_com_n_241, A2 => fsm_com_n_24, B => fsm_com_n_274, Z => fsm_com_n_289);
  fsm_com_g21121 : OAI211D1BWP7T port map(A1 => fsm_com_n_164, A2 => fsm_com_n_536, B => fsm_com_n_550, C => fsm_com_energy(3), ZN => fsm_com_n_288);
  fsm_com_g21122 : OAI21D0BWP7T port map(A1 => fsm_com_n_48, A2 => FE_PHN383_energy_d_10, B => fsm_com_n_253, ZN => fsm_com_n_297);
  fsm_com_g21123 : AOI221D0BWP7T port map(A1 => fsm_com_n_550, A2 => fsm_com_n_77, B1 => fsm_com_n_549, B2 => fsm_com_n_51, C => fsm_com_n_269, ZN => fsm_com_n_296);
  fsm_com_g21124 : NR2XD0BWP7T port map(A1 => fsm_com_n_268, A2 => fsm_com_energy(6), ZN => fsm_com_n_295);
  fsm_com_g21125 : NR2XD0BWP7T port map(A1 => fsm_com_n_266, A2 => yplayer(0), ZN => fsm_com_n_294);
  fsm_com_g21130 : OAI21D0BWP7T port map(A1 => fsm_com_n_234, A2 => fsm_com_n_50, B => fsm_com_n_550, ZN => fsm_com_n_281);
  fsm_com_g21133 : AOI211XD0BWP7T port map(A1 => fsm_com_n_122, A2 => xplayer(2), B => fsm_com_n_247, C => fsm_com_n_127, ZN => fsm_com_n_278);
  fsm_com_g21134 : MAOI22D0BWP7T port map(A1 => fsm_com_n_246, A2 => fsm_com_energy(4), B1 => fsm_com_n_118, B2 => FE_PHN224_fsm_com_reached_high_0, ZN => fsm_com_n_277);
  fsm_com_g21135 : AO21D0BWP7T port map(A1 => fsm_com_n_549, A2 => FE_PHN233_fsm_com_n_22, B => fsm_com_n_269, Z => fsm_com_n_276);
  fsm_com_g21136 : OA21D0BWP7T port map(A1 => fsm_com_n_181, A2 => fsm_com_n_96, B => fsm_com_n_255, Z => fsm_com_n_275);
  fsm_com_g21137 : ND3D0BWP7T port map(A1 => fsm_com_n_245, A2 => fsm_com_n_141, A3 => fsm_com_n_538, ZN => fsm_com_n_286);
  fsm_com_g21138 : AO21D0BWP7T port map(A1 => fsm_com_n_185, A2 => fsm_com_n_100, B => fsm_com_n_259, Z => fsm_com_n_285);
  fsm_com_g21139 : OAI21D0BWP7T port map(A1 => fsm_com_n_182, A2 => fsm_com_n_99, B => fsm_com_n_254, ZN => fsm_com_n_284);
  fsm_com_g21140 : OAI21D0BWP7T port map(A1 => fsm_com_n_74, A2 => energy_d(6), B => fsm_com_n_262, ZN => fsm_com_n_283);
  fsm_com_g21141 : AOI22D0BWP7T port map(A1 => fsm_com_n_140, A2 => fsm_com_n_14, B1 => FE_PHN224_fsm_com_reached_high_0, B2 => fsm_com_reached_high(1), ZN => fsm_com_n_282);
  fsm_com_g21142 : CKND1BWP7T port map(I => fsm_com_n_271, ZN => fsm_com_n_272);
  fsm_com_g21143 : INVD1BWP7T port map(I => fsm_com_n_264, ZN => fsm_com_n_265);
  fsm_com_g21144 : ND3D0BWP7T port map(A1 => fsm_com_n_201, A2 => fsm_com_n_538, A3 => FE_DBTN0_reset, ZN => fsm_com_n_263);
  fsm_com_g21145 : ND2D1BWP7T port map(A1 => fsm_com_n_241, A2 => fsm_com_n_24, ZN => fsm_com_n_274);
  fsm_com_g21146 : AOI21D0BWP7T port map(A1 => fsm_com_n_203, A2 => fsm_com_n_24, B => fsm_com_n_70, ZN => fsm_com_n_273);
  fsm_com_g21147 : ND2D1BWP7T port map(A1 => fsm_com_n_230, A2 => fsm_com_n_30, ZN => fsm_com_n_271);
  fsm_com_g21148 : IND2D1BWP7T port map(A1 => fsm_com_n_568, B1 => fsm_com_n_230, ZN => fsm_com_n_270);
  fsm_com_g21149 : IND3D1BWP7T port map(A1 => fsm_com_n_55, B1 => fsm_com_n_75, B2 => fsm_com_n_213, ZN => fsm_com_n_269);
  fsm_com_g21150 : ND2D1BWP7T port map(A1 => fsm_com_n_241, A2 => fsm_com_n_84, ZN => fsm_com_n_268);
  fsm_com_g21152 : ND2D1BWP7T port map(A1 => fsm_com_n_230, A2 => fsm_com_n_568, ZN => fsm_com_n_266);
  fsm_com_g21153 : IAO21D0BWP7T port map(A1 => fsm_com_n_203, A2 => fsm_com_n_70, B => fsm_com_n_189, ZN => fsm_com_n_264);
  fsm_com_g21156 : INVD0BWP7T port map(I => fsm_com_n_257, ZN => fsm_com_n_258);
  fsm_com_g21157 : MAOI22D0BWP7T port map(A1 => fsm_com_n_172, A2 => yplayer(3), B1 => fsm_com_n_172, B2 => yplayer(3), ZN => fsm_com_n_251);
  fsm_com_g21158 : OA21D0BWP7T port map(A1 => fsm_com_n_205, A2 => fsm_com_n_180, B => fsm_com_n_69, Z => fsm_com_n_250);
  fsm_com_g21159 : MOAI22D0BWP7T port map(A1 => fsm_com_n_167, A2 => FE_PHN232_energy_d_7, B1 => fsm_com_n_167, B2 => FE_PHN232_energy_d_7, ZN => fsm_com_n_262);
  fsm_com_g21160 : OR3D1BWP7T port map(A1 => fsm_com_n_194, A2 => fsm_com_n_242, A3 => fsm_com_n_139, Z => fsm_com_n_261);
  fsm_com_g21161 : MOAI22D0BWP7T port map(A1 => fsm_com_n_169, A2 => energy_d(3), B1 => fsm_com_n_169, B2 => energy_d(3), ZN => fsm_com_n_260);
  fsm_com_g21162 : MAOI22D0BWP7T port map(A1 => fsm_com_n_175, A2 => level_d(3), B1 => fsm_com_n_175, B2 => level_d(3), ZN => fsm_com_n_259);
  fsm_com_g21163 : AOI21D0BWP7T port map(A1 => fsm_com_n_95, A2 => fsm_com_n_186, B => fsm_com_n_54, ZN => fsm_com_n_257);
  fsm_com_g21164 : MOAI22D0BWP7T port map(A1 => fsm_com_n_174, A2 => level_d(7), B1 => fsm_com_n_174, B2 => level_d(7), ZN => fsm_com_n_256);
  fsm_com_g21165 : MOAI22D0BWP7T port map(A1 => fsm_com_n_173, A2 => score_d(15), B1 => fsm_com_n_173, B2 => score_d(15), ZN => fsm_com_n_255);
  fsm_com_g21166 : MOAI22D0BWP7T port map(A1 => fsm_com_n_170, A2 => score_d(11), B1 => fsm_com_n_170, B2 => score_d(11), ZN => fsm_com_n_254);
  fsm_com_g21167 : MOAI22D0BWP7T port map(A1 => fsm_com_n_165, A2 => energy_d(11), B1 => fsm_com_n_165, B2 => energy_d(11), ZN => fsm_com_n_253);
  fsm_com_g21168 : AO21D0BWP7T port map(A1 => fsm_com_n_168, A2 => fsm_com_energy(3), B => fsm_com_n_243, Z => fsm_com_n_252);
  fsm_com_g21169 : INVD0BWP7T port map(I => fsm_com_n_241, ZN => fsm_com_n_240);
  fsm_com_g21170 : CKND2D0BWP7T port map(A1 => fsm_com_n_210, A2 => fsm_com_energy(5), ZN => fsm_com_n_238);
  fsm_com_g21171 : CKND2D0BWP7T port map(A1 => fsm_com_n_210, A2 => fsm_com_energy(7), ZN => fsm_com_n_237);
  fsm_com_g21172 : CKND2D0BWP7T port map(A1 => fsm_com_n_210, A2 => fsm_com_energy(6), ZN => fsm_com_n_236);
  fsm_com_g21173 : INR2D0BWP7T port map(A1 => fsm_com_energy(3), B1 => fsm_com_n_209, ZN => fsm_com_n_235);
  fsm_com_g21174 : ND2D1BWP7T port map(A1 => fsm_com_n_203, A2 => fsm_com_n_4, ZN => fsm_com_n_249);
  fsm_com_g21175 : INR2D0BWP7T port map(A1 => fsm_com_n_180, B1 => fsm_com_n_209, ZN => fsm_com_n_248);
  fsm_com_g21176 : NR2D0BWP7T port map(A1 => fsm_com_n_213, A2 => fsm_com_n_35, ZN => fsm_com_n_247);
  fsm_com_g21177 : OR2D1BWP7T port map(A1 => fsm_com_n_139, A2 => fsm_com_n_219, Z => fsm_com_n_246);
  fsm_com_g21178 : NR4D0BWP7T port map(A1 => fsm_com_n_163, A2 => fsm_com_n_550, A3 => fsm_com_n_547, A4 => fsm_com_n_66, ZN => fsm_com_n_245);
  fsm_com_g21179 : NR2D0BWP7T port map(A1 => fsm_com_n_209, A2 => fsm_com_n_4, ZN => fsm_com_n_244);
  fsm_com_g21180 : NR2XD0BWP7T port map(A1 => fsm_com_n_168, A2 => fsm_com_energy(3), ZN => fsm_com_n_243);
  fsm_com_g21181 : AN2D1BWP7T port map(A1 => fsm_com_n_205, A2 => fsm_com_n_69, Z => fsm_com_n_242);
  fsm_com_g21182 : NR2XD0BWP7T port map(A1 => fsm_com_n_164, A2 => fsm_com_energy(3), ZN => fsm_com_n_241);
  fsm_com_g21183 : NR2D1BWP7T port map(A1 => fsm_com_n_209, A2 => fsm_com_n_212, ZN => fsm_com_n_239);
  fsm_com_g21184 : INVD1BWP7T port map(I => fsm_com_n_602, ZN => fsm_com_n_228);
  fsm_com_g21185 : MAOI22D0BWP7T port map(A1 => fsm_com_n_193, A2 => FE_PHN188_fsm_com_n_28, B1 => fsm_com_n_193, B2 => FE_PHN188_fsm_com_n_28, ZN => fsm_com_n_227);
  fsm_com_g21186 : OR2D1BWP7T port map(A1 => fsm_com_n_184, A2 => fsm_com_n_98, Z => fsm_com_n_226);
  fsm_com_g21187 : MOAI22D0BWP7T port map(A1 => fsm_com_n_65, A2 => fsm_com_n_150, B1 => fsm_com_n_137, B2 => level_abs(3), ZN => fsm_com_n_225);
  fsm_com_g21188 : OAI22D0BWP7T port map(A1 => fsm_com_n_189, A2 => fsm_com_energy(1), B1 => fsm_com_n_557, B2 => fsm_com_n_536, ZN => fsm_com_n_224);
  fsm_com_g21189 : MAOI22D0BWP7T port map(A1 => fsm_com_n_140, A2 => level_abs(4), B1 => fsm_com_n_140, B2 => level_abs(4), ZN => fsm_com_n_223);
  fsm_com_g21190 : OAI211D1BWP7T port map(A1 => fsm_com_n_160, A2 => fsm_com_n_117, B => fsm_com_n_101, C => fsm_com_n_603, ZN => fsm_com_n_222);
  fsm_com_g21191 : OAI211D1BWP7T port map(A1 => fsm_com_n_31, A2 => fsm_com_n_153, B => fsm_com_n_188, C => fsm_com_n_195, ZN => fsm_com_n_221);
  fsm_com_g21192 : OAI211D1BWP7T port map(A1 => fsm_com_n_159, A2 => fsm_com_n_117, B => fsm_com_n_90, C => fsm_com_n_604, ZN => fsm_com_n_220);
  fsm_com_g21193 : OAI21D0BWP7T port map(A1 => fsm_com_n_536, A2 => fsm_com_n_77, B => fsm_com_n_213, ZN => fsm_com_n_234);
  fsm_com_g21194 : INR2D1BWP7T port map(A1 => fsm_com_n_217, B1 => fsm_com_n_218, ZN => fsm_com_n_233);
  fsm_com_g21195 : AOI221D0BWP7T port map(A1 => fsm_com_n_146, A2 => level_abs(2), B1 => fsm_com_n_133, B2 => fsm_com_n_25, C => FE_PHN224_fsm_com_reached_high_0, ZN => fsm_com_n_232);
  fsm_com_g21196 : MOAI22D0BWP7T port map(A1 => fsm_com_n_190, A2 => fsm_com_n_5, B1 => fsm_com_n_190, B2 => fsm_com_n_5, ZN => fsm_com_n_231);
  fsm_com_g21197 : NR3D0BWP7T port map(A1 => fsm_com_n_1, A2 => fsm_com_n_549, A3 => fsm_com_n_550, ZN => fsm_com_n_230);
  fsm_com_g21199 : INVD0BWP7T port map(I => fsm_com_n_212, ZN => fsm_com_n_211);
  fsm_com_g21200 : INVD1BWP7T port map(I => fsm_com_n_210, ZN => fsm_com_n_209);
  fsm_com_g21201 : IND3D0BWP7T port map(A1 => fsm_com_n_0, B1 => animation_done, B2 => fsm_com_n_545, ZN => fsm_com_n_208);
  fsm_com_g21202 : IND2D1BWP7T port map(A1 => fsm_com_n_194, B1 => fsm_com_n_75, ZN => fsm_com_n_219);
  fsm_com_g21203 : INR2D1BWP7T port map(A1 => fsm_com_n_196, B1 => score_d(1), ZN => fsm_com_n_218);
  fsm_com_g21204 : IND2D1BWP7T port map(A1 => fsm_com_n_196, B1 => score_d(1), ZN => fsm_com_n_217);
  fsm_com_g21205 : ND2D1BWP7T port map(A1 => fsm_com_n_193, A2 => score_d(0), ZN => fsm_com_n_216);
  fsm_com_g21206 : NR2XD0BWP7T port map(A1 => fsm_com_n_190, A2 => energy_d(0), ZN => fsm_com_n_215);
  fsm_com_g21207 : IND2D1BWP7T port map(A1 => fsm_com_n_192, B1 => fsm_com_n_545, ZN => fsm_com_n_214);
  fsm_com_g21208 : INR2XD0BWP7T port map(A1 => fsm_com_n_58, B1 => fsm_com_n_1, ZN => fsm_com_n_213);
  fsm_com_g21209 : INR2XD0BWP7T port map(A1 => fsm_com_n_191, B1 => fsm_com_n_539, ZN => fsm_com_n_212);
  fsm_com_g21210 : IND2D1BWP7T port map(A1 => fsm_com_n_559, B1 => fsm_com_n_191, ZN => fsm_com_n_210);
  fsm_com_g21211 : OAI32D1BWP7T port map(A1 => level_abs(1), A2 => fsm_com_n_16, A3 => fsm_com_n_65, B1 => fsm_com_n_21, B2 => fsm_com_n_161, ZN => fsm_com_n_202);
  fsm_com_g21212 : AOI211XD0BWP7T port map(A1 => fsm_com_n_137, A2 => level_abs(0), B => fsm_com_n_124, C => fsm_com_n_544, ZN => fsm_com_n_201);
  fsm_com_g21213 : NR3D0BWP7T port map(A1 => fsm_com_n_155, A2 => fsm_com_n_550, A3 => fsm_com_n_91, ZN => fsm_com_n_200);
  fsm_com_g21214 : AO21D0BWP7T port map(A1 => fsm_com_n_153, A2 => fsm_com_n_555, B => fsm_com_n_194, Z => fsm_com_n_199);
  fsm_com_g21215 : OAI32D1BWP7T port map(A1 => fsm_com_energy(1), A2 => fsm_com_n_91, A3 => fsm_com_n_68, B1 => fsm_com_n_557, B2 => fsm_com_n_550, ZN => fsm_com_n_198);
  fsm_com_g21216 : OAI22D0BWP7T port map(A1 => fsm_com_n_161, A2 => fsm_com_n_25, B1 => fsm_com_n_65, B2 => fsm_com_n_125, ZN => FE_PHN356_fsm_com_n_197);
  fsm_com_g21217 : OAI22D0BWP7T port map(A1 => fsm_com_n_156, A2 => fsm_com_n_555, B1 => fsm_com_n_154, B2 => fsm_com_n_557, ZN => fsm_com_n_207);
  fsm_com_g21218 : OAI22D0BWP7T port map(A1 => fsm_com_n_155, A2 => fsm_com_n_555, B1 => fsm_com_n_153, B2 => fsm_com_n_557, ZN => fsm_com_n_206);
  fsm_com_g21219 : MAOI22D0BWP7T port map(A1 => fsm_com_n_157, A2 => fsm_com_n_31, B1 => fsm_com_n_153, B2 => fsm_com_n_561, ZN => fsm_com_n_205);
  fsm_com_g21220 : OAI21D0BWP7T port map(A1 => fsm_com_n_157, A2 => fsm_com_n_32, B => fsm_com_n_75, ZN => fsm_com_n_204);
  fsm_com_g21221 : OAI22D0BWP7T port map(A1 => fsm_com_n_154, A2 => fsm_com_n_561, B1 => fsm_com_n_157, B2 => fsm_com_n_555, ZN => fsm_com_n_203);
  fsm_com_g21222 : INVD1BWP7T port map(I => fsm_com_n_188, ZN => fsm_com_n_189);
  fsm_com_g21223 : AOI22D0BWP7T port map(A1 => fsm_com_n_135, A2 => fsm_com_n_144, B1 => fsm_com_n_121, B2 => fsm_com_energy(1), ZN => fsm_com_n_187);
  fsm_com_g21225 : AOI221D0BWP7T port map(A1 => fsm_com_n_559, A2 => fsm_com_n_107, B1 => fsm_com_n_561, B2 => fsm_com_n_39, C => fsm_com_n_128, ZN => fsm_com_n_196);
  fsm_com_g21226 : ND2D1BWP7T port map(A1 => fsm_com_n_157, A2 => fsm_com_n_561, ZN => fsm_com_n_195);
  fsm_com_g21227 : NR2D1BWP7T port map(A1 => fsm_com_n_156, A2 => fsm_com_n_36, ZN => fsm_com_n_194);
  fsm_com_g21228 : OAI211D1BWP7T port map(A1 => fsm_com_n_110, A2 => fsm_com_n_32, B => fsm_com_n_148, C => fsm_com_n_129, ZN => fsm_com_n_193);
  fsm_com_g21229 : OAI21D0BWP7T port map(A1 => fsm_com_n_133, A2 => fsm_com_n_25, B => fsm_com_n_147, ZN => fsm_com_n_192);
  fsm_com_g21230 : NR2XD0BWP7T port map(A1 => fsm_com_n_171, A2 => fsm_com_n_37, ZN => fsm_com_n_191);
  fsm_com_g21231 : INR3D0BWP7T port map(A1 => fsm_com_n_158, B1 => dir_mined(1), B2 => fsm_com_n_558, ZN => fsm_com_n_190);
  fsm_com_g21232 : ND2D1BWP7T port map(A1 => fsm_com_n_156, A2 => fsm_com_n_557, ZN => fsm_com_n_188);
  fsm_com_g21233 : MAOI22D0BWP7T port map(A1 => fsm_com_n_79, A2 => yplayer(2), B1 => fsm_com_n_79, B2 => yplayer(2), ZN => fsm_com_n_179);
  fsm_com_g21234 : OAI21D0BWP7T port map(A1 => fsm_com_n_74, A2 => fsm_com_n_18, B => fsm_com_n_167, ZN => fsm_com_n_178);
  fsm_com_g21235 : OA21D0BWP7T port map(A1 => fsm_com_n_48, A2 => fsm_com_n_19, B => fsm_com_n_165, Z => fsm_com_n_177);
  fsm_com_g21236 : MAOI22D0BWP7T port map(A1 => fsm_com_n_42, A2 => xplayer(1), B1 => fsm_com_n_44, B2 => fsm_com_n_89, ZN => fsm_com_n_176);
  fsm_com_g21237 : OA21D0BWP7T port map(A1 => fsm_com_n_62, A2 => fsm_com_n_15, B => fsm_com_n_164, Z => fsm_com_n_186);
  fsm_com_g21238 : MAOI22D0BWP7T port map(A1 => fsm_com_n_57, A2 => level_d(2), B1 => fsm_com_n_57, B2 => level_d(2), ZN => fsm_com_n_185);
  fsm_com_g21239 : MOAI22D0BWP7T port map(A1 => fsm_com_n_56, A2 => level_d(6), B1 => fsm_com_n_56, B2 => level_d(6), ZN => fsm_com_n_184);
  fsm_com_g21240 : MAOI22D0BWP7T port map(A1 => fsm_com_n_47, A2 => fsm_com_n_13, B1 => fsm_com_n_47, B2 => fsm_com_n_13, ZN => fsm_com_n_183);
  fsm_com_g21241 : MOAI22D0BWP7T port map(A1 => fsm_com_n_49, A2 => score_d(10), B1 => fsm_com_n_49, B2 => score_d(10), ZN => fsm_com_n_182);
  fsm_com_g21242 : MOAI22D0BWP7T port map(A1 => fsm_com_n_76, A2 => score_d(14), B1 => fsm_com_n_76, B2 => score_d(14), ZN => fsm_com_n_181);
  fsm_com_g21243 : OAI21D0BWP7T port map(A1 => fsm_com_n_86, A2 => fsm_com_n_15, B => fsm_com_n_168, ZN => fsm_com_n_180);
  fsm_com_g21245 : ND2D0BWP7T port map(A1 => fsm_com_n_132, A2 => fsm_com_n_54, ZN => fsm_com_n_163);
  fsm_com_g21246 : NR2XD0BWP7T port map(A1 => fsm_com_n_142, A2 => button_left, ZN => fsm_com_n_162);
  fsm_com_g21247 : IND2D1BWP7T port map(A1 => fsm_com_n_57, B1 => level_d(2), ZN => fsm_com_n_175);
  fsm_com_g21248 : IND2D1BWP7T port map(A1 => fsm_com_n_56, B1 => level_d(6), ZN => fsm_com_n_174);
  fsm_com_g21249 : IND2D1BWP7T port map(A1 => fsm_com_n_76, B1 => score_d(14), ZN => fsm_com_n_173);
  fsm_com_g21250 : OR2D1BWP7T port map(A1 => fsm_com_n_79, A2 => fsm_com_n_10, Z => fsm_com_n_172);
  fsm_com_g21251 : IND2D1BWP7T port map(A1 => fsm_com_n_546, B1 => fsm_com_n_141, ZN => fsm_com_n_171);
  fsm_com_g21252 : IND2D1BWP7T port map(A1 => fsm_com_n_49, B1 => score_d(10), ZN => fsm_com_n_170);
  fsm_com_g21253 : AN2D0BWP7T port map(A1 => fsm_com_n_47, A2 => energy_d(2), Z => fsm_com_n_169);
  fsm_com_g21254 : ND2D1BWP7T port map(A1 => fsm_com_n_86, A2 => fsm_com_n_15, ZN => fsm_com_n_168);
  fsm_com_g21255 : ND2D1BWP7T port map(A1 => fsm_com_n_74, A2 => fsm_com_n_18, ZN => fsm_com_n_167);
  fsm_com_g21256 : ND2D1BWP7T port map(A1 => fsm_com_n_126, A2 => score_d(7), ZN => fsm_com_n_166);
  fsm_com_g21257 : ND2D1BWP7T port map(A1 => fsm_com_n_48, A2 => fsm_com_n_19, ZN => fsm_com_n_165);
  fsm_com_g21258 : ND2D1BWP7T port map(A1 => fsm_com_n_62, A2 => fsm_com_n_15, ZN => fsm_com_n_164);
  fsm_com_g21259 : CKND1BWP7T port map(I => fsm_com_n_159, ZN => fsm_com_n_160);
  fsm_com_g21260 : INVD0BWP7T port map(I => fsm_com_n_156, ZN => fsm_com_n_155);
  fsm_com_g21261 : INVD1BWP7T port map(I => fsm_com_n_154, ZN => fsm_com_n_153);
  fsm_com_g21262 : INVD1BWP7T port map(I => fsm_com_n_152, ZN => fsm_com_n_151);
  fsm_com_g21263 : MAOI22D0BWP7T port map(A1 => fsm_com_n_120, A2 => level_abs(3), B1 => fsm_com_n_120, B2 => level_abs(3), ZN => fsm_com_n_150);
  fsm_com_g21265 : AOI33D1BWP7T port map(A1 => fsm_com_n_557, A2 => fsm_com_n_60, A3 => map_data(37), B1 => fsm_com_n_555, B2 => fsm_com_n_87, B3 => map_data(34), ZN => fsm_com_n_148);
  fsm_com_g21266 : ND4D0BWP7T port map(A1 => fsm_com_n_52, A2 => fsm_com_n_78, A3 => level_abs(1), A4 => level_abs(3), ZN => fsm_com_n_147);
  fsm_com_g21267 : AO211D0BWP7T port map(A1 => fsm_com_n_78, A2 => fsm_com_n_21, B => fsm_com_n_53, C => level_abs(3), Z => fsm_com_n_146);
  fsm_com_g21268 : NR3D0BWP7T port map(A1 => fsm_com_n_117, A2 => fsm_com_n_59, A3 => button_left, ZN => fsm_com_n_145);
  fsm_com_g21269 : NR2D1BWP7T port map(A1 => fsm_com_n_137, A2 => fsm_com_n_124, ZN => fsm_com_n_161);
  fsm_com_g21270 : IOA21D1BWP7T port map(A1 => button_left, A2 => button_mining, B => fsm_com_n_142, ZN => fsm_com_n_159);
  fsm_com_g21272 : NR2XD0BWP7T port map(A1 => fsm_com_n_138, A2 => fsm_com_n_68, ZN => fsm_com_n_158);
  fsm_com_g21273 : AOI221D0BWP7T port map(A1 => fsm_com_n_63, A2 => map_data(19), B1 => map_data(18), B2 => map_data(20), C => fsm_com_n_571, ZN => fsm_com_n_157);
  fsm_com_g21274 : AOI221D0BWP7T port map(A1 => fsm_com_n_61, A2 => map_data(37), B1 => map_data(36), B2 => map_data(38), C => fsm_com_n_565, ZN => fsm_com_n_156);
  fsm_com_g21275 : AOI221D0BWP7T port map(A1 => fsm_com_n_88, A2 => map_data(34), B1 => map_data(33), B2 => map_data(35), C => fsm_com_n_568, ZN => fsm_com_n_154);
  fsm_com_g21276 : NR2XD0BWP7T port map(A1 => fsm_com_n_136, A2 => FE_OFN0_reset, ZN => fsm_com_n_152);
  fsm_com_g21277 : INVD0BWP7T port map(I => fsm_com_n_91, ZN => fsm_com_n_144);
  fsm_com_g21278 : INVD1BWP7T port map(I => fsm_com_n_136, ZN => fsm_com_n_137);
  fsm_com_g21279 : ND2D1BWP7T port map(A1 => fsm_com_n_119, A2 => fsm_com_n_4, ZN => fsm_com_n_135);
  fsm_com_g21281 : IAO21D0BWP7T port map(A1 => fsm_com_n_65, A2 => FE_PHN205_fsm_com_reached_high_1, B => fsm_com_n_544, ZN => fsm_com_n_143);
  fsm_com_g21282 : OAI21D0BWP7T port map(A1 => fsm_com_n_38, A2 => button_right, B => button_mining, ZN => fsm_com_n_142);
  fsm_com_g21283 : NR3D0BWP7T port map(A1 => fsm_com_n_82, A2 => fsm_com_n_46, A3 => fsm_com_n_85, ZN => fsm_com_n_141);
  fsm_com_g21284 : IND2D1BWP7T port map(A1 => fsm_com_n_120, B1 => level_abs(3), ZN => fsm_com_n_140);
  fsm_com_g21285 : OR2D1BWP7T port map(A1 => fsm_com_n_121, A2 => fsm_com_n_55, Z => fsm_com_n_139);
  fsm_com_g21286 : ND2D1BWP7T port map(A1 => fsm_com_n_119, A2 => fsm_com_n_73, ZN => fsm_com_n_138);
  fsm_com_g21287 : ND3D0BWP7T port map(A1 => fsm_com_n_83, A2 => fsm_com_n_65, A3 => fsm_com_n_538, ZN => fsm_com_n_136);
  fsm_com_g21288 : MAOI22D0BWP7T port map(A1 => fsm_com_n_42, A2 => xplayer(0), B1 => fsm_com_n_44, B2 => yplayer(0), ZN => fsm_com_n_131);
  fsm_com_g21289 : AOI21D0BWP7T port map(A1 => fsm_com_n_67, A2 => fsm_com_n_73, B => xplayer(0), ZN => fsm_com_n_130);
  fsm_com_g21290 : IIND4D0BWP7T port map(A1 => map_data(51), A2 => map_data(53), B1 => fsm_com_n_559, B2 => map_data(52), ZN => fsm_com_n_129);
  fsm_com_g21291 : OAI33D1BWP7T port map(A1 => map_data(36), A2 => fsm_com_n_566, A3 => fsm_com_n_36, B1 => map_data(33), B2 => fsm_com_n_569, B3 => fsm_com_n_31, ZN => fsm_com_n_128);
  fsm_com_g21292 : NR3D0BWP7T port map(A1 => fsm_com_n_67, A2 => fsm_com_n_77, A3 => xplayer(2), ZN => fsm_com_n_127);
  fsm_com_g21293 : AOI31D0BWP7T port map(A1 => FE_PHN244_score_d_4, A2 => score_d(6), A3 => score_d(5), B => fsm_com_n_108, ZN => fsm_com_n_126);
  fsm_com_g21294 : AOI32D1BWP7T port map(A1 => fsm_com_n_25, A2 => level_abs(1), A3 => level_abs(0), B1 => fsm_com_n_21, B2 => level_abs(2), ZN => fsm_com_n_125);
  fsm_com_g21295 : ND3D0BWP7T port map(A1 => fsm_com_n_52, A2 => fsm_com_n_21, A3 => level_abs(3), ZN => fsm_com_n_133);
  fsm_com_g21296 : NR3D0BWP7T port map(A1 => fsm_com_n_81, A2 => fsm_com_n_559, A3 => fsm_com_n_561, ZN => fsm_com_n_132);
  fsm_com_g21297 : INVD1BWP7T port map(I => fsm_com_n_115, ZN => fsm_com_n_114);
  fsm_com_g21298 : AO21D0BWP7T port map(A1 => energy_d(5), A2 => energy_d(4), B => fsm_com_n_74, Z => fsm_com_n_113);
  fsm_com_g21299 : AOI21D0BWP7T port map(A1 => energy_d(9), A2 => energy_d(8), B => fsm_com_n_48, ZN => fsm_com_n_112);
  fsm_com_g21300 : ND2D1BWP7T port map(A1 => fsm_com_n_71, A2 => energy_d(0), ZN => fsm_com_n_111);
  fsm_com_g21301 : IND2D1BWP7T port map(A1 => fsm_com_n_63, B1 => map_data(19), ZN => fsm_com_n_110);
  fsm_com_g21303 : NR3D0BWP7T port map(A1 => score_d(5), A2 => FE_PHN244_score_d_4, A3 => score_d(6), ZN => fsm_com_n_108);
  fsm_com_g21304 : INR3D0BWP7T port map(A1 => map_data(53), B1 => map_data(51), B2 => map_data(52), ZN => fsm_com_n_107);
  fsm_com_g21305 : NR2XD0BWP7T port map(A1 => fsm_com_n_65, A2 => level_abs(0), ZN => fsm_com_n_124);
  fsm_com_g21306 : CKAN2D1BWP7T port map(A1 => fsm_com_n_67, A2 => fsm_com_n_44, Z => fsm_com_n_123);
  fsm_com_g21307 : NR2XD0BWP7T port map(A1 => fsm_com_n_73, A2 => fsm_com_n_51, ZN => fsm_com_n_122);
  fsm_com_g21308 : OAI21D0BWP7T port map(A1 => fsm_com_n_30, A2 => fsm_com_n_568, B => fsm_com_n_41, ZN => fsm_com_n_121);
  fsm_com_g21309 : OR2D1BWP7T port map(A1 => fsm_com_n_78, A2 => fsm_com_n_21, Z => fsm_com_n_120);
  fsm_com_g21310 : AOI21D0BWP7T port map(A1 => fsm_com_n_548, A2 => fsm_com_n_568, B => fsm_com_n_43, ZN => fsm_com_n_119);
  fsm_com_g21311 : ND2D1BWP7T port map(A1 => fsm_com_n_66, A2 => FE_PHN205_fsm_com_reached_high_1, ZN => fsm_com_n_118);
  fsm_com_g21312 : ND2D1BWP7T port map(A1 => fsm_com_n_82, A2 => vga_done, ZN => fsm_com_n_117);
  fsm_com_g21313 : ND2D1BWP7T port map(A1 => fsm_com_n_66, A2 => FE_PHN224_fsm_com_reached_high_0, ZN => fsm_com_n_116);
  fsm_com_g21314 : ND2D1BWP7T port map(A1 => fsm_com_n_66, A2 => FE_DBTN0_reset, ZN => fsm_com_n_115);
  fsm_com_g21315 : INVD0BWP7T port map(I => fsm_com_n_92, ZN => fsm_com_n_93);
  fsm_com_g21316 : AOI22D0BWP7T port map(A1 => fsm_com_n_549, A2 => fsm_com_n_570, B1 => fsm_com_n_547, B2 => fsm_com_n_564, ZN => fsm_com_n_90);
  fsm_com_g21317 : AOI22D0BWP7T port map(A1 => fsm_com_n_8, A2 => yplayer(0), B1 => fsm_com_n_11, B2 => yplayer(1), ZN => fsm_com_n_89);
  fsm_com_g21318 : AOI22D0BWP7T port map(A1 => fsm_com_n_7, A2 => energy_d(0), B1 => fsm_com_n_5, B2 => FE_PHN403_energy_d_1, ZN => fsm_com_n_106);
  fsm_com_g21319 : IND4D0BWP7T port map(A1 => fsm_com_edge_detec3(2), B1 => fsm_com_edge_detec2(2), B2 => fsm_com_edge_detec1(2), B3 => fsm_com_edge_detec0(2), ZN => fsm_com_n_105);
  fsm_com_g21320 : OAI22D0BWP7T port map(A1 => fsm_com_n_29, A2 => fsm_com_n_570, B1 => fsm_com_n_33, B2 => fsm_com_n_564, ZN => fsm_com_n_104);
  fsm_com_g21321 : IND4D0BWP7T port map(A1 => fsm_com_edge_detec3(3), B1 => FE_PHN212_fsm_com_edge_detec2_3, B2 => fsm_com_edge_detec1(3), B3 => FE_PHN209_fsm_com_edge_detec0_3, ZN => fsm_com_n_103);
  fsm_com_g21322 : OAI22D0BWP7T port map(A1 => fsm_com_n_549, A2 => fsm_com_n_568, B1 => fsm_com_n_548, B2 => fsm_com_n_571, ZN => fsm_com_n_102);
  fsm_com_g21323 : MAOI22D0BWP7T port map(A1 => fsm_com_n_550, A2 => fsm_com_n_537, B1 => fsm_com_n_30, B2 => fsm_com_n_567, ZN => fsm_com_n_101);
  fsm_com_g21324 : XNR2D1BWP7T port map(A1 => level_d(0), A2 => FE_PHN454_level_d_1, ZN => fsm_com_n_100);
  fsm_com_g21325 : CKXOR2D1BWP7T port map(A1 => FE_PHN249_score_d_8, A2 => score_d(9), Z => fsm_com_n_99);
  fsm_com_g21326 : CKXOR2D1BWP7T port map(A1 => level_d(4), A2 => level_d(5), Z => fsm_com_n_98);
  fsm_com_g21327 : MOAI22D0BWP7T port map(A1 => dir_mined(2), A2 => FE_PHN403_energy_d_1, B1 => dir_mined(2), B2 => FE_PHN403_energy_d_1, ZN => fsm_com_n_97);
  fsm_com_g21328 : CKXOR2D1BWP7T port map(A1 => FE_PHN227_score_d_12, A2 => score_d(13), Z => fsm_com_n_96);
  fsm_com_g21329 : AO22D0BWP7T port map(A1 => fsm_com_n_30, A2 => fsm_com_n_571, B1 => fsm_com_n_568, B2 => fsm_com_n_29, Z => fsm_com_n_95);
  fsm_com_g21330 : IND4D0BWP7T port map(A1 => fsm_com_edge_detec3(0), B1 => fsm_com_edge_detec2(0), B2 => fsm_com_edge_detec1(0), B3 => fsm_com_edge_detec0(0), ZN => fsm_com_n_94);
  fsm_com_g21331 : IND4D0BWP7T port map(A1 => fsm_com_edge_detec3(1), B1 => fsm_com_edge_detec2(1), B2 => fsm_com_edge_detec1(1), B3 => fsm_com_edge_detec0(1), ZN => fsm_com_n_92);
  fsm_com_g21332 : MOAI22D0BWP7T port map(A1 => fsm_com_n_4, A2 => fsm_com_energy(0), B1 => fsm_com_n_4, B2 => fsm_com_energy(0), ZN => fsm_com_n_91);
  fsm_com_g21333 : CKND1BWP7T port map(I => fsm_com_n_87, ZN => fsm_com_n_88);
  fsm_com_g21334 : INVD0BWP7T port map(I => fsm_com_n_81, ZN => fsm_com_n_80);
  fsm_com_g21335 : INVD0BWP7T port map(I => fsm_com_n_73, ZN => fsm_com_n_72);
  fsm_com_g21336 : INVD1BWP7T port map(I => fsm_com_n_70, ZN => fsm_com_n_69);
  fsm_com_g21337 : INVD1BWP7T port map(I => fsm_com_n_68, ZN => fsm_com_n_67);
  fsm_com_g21338 : INVD1BWP7T port map(I => fsm_com_n_66, ZN => fsm_com_n_65);
  fsm_com_g21339 : NR2XD0BWP7T port map(A1 => fsm_com_n_568, A2 => xplayer(0), ZN => fsm_com_n_64);
  fsm_com_g21340 : NR2D1BWP7T port map(A1 => map_data(35), A2 => map_data(33), ZN => fsm_com_n_87);
  fsm_com_g21341 : CKND2D1BWP7T port map(A1 => fsm_com_energy(0), A2 => fsm_com_energy(1), ZN => fsm_com_n_86);
  fsm_com_g21342 : NR2D1BWP7T port map(A1 => fsm_com_n_563, A2 => fsm_com_n_556, ZN => fsm_com_n_85);
  fsm_com_g21343 : NR2XD0BWP7T port map(A1 => fsm_com_energy(4), A2 => fsm_com_energy(5), ZN => fsm_com_n_84);
  fsm_com_g21344 : NR2XD0BWP7T port map(A1 => fsm_com_n_545, A2 => fsm_com_n_544, ZN => fsm_com_n_83);
  fsm_com_g21345 : NR2D0BWP7T port map(A1 => fsm_com_n_551, A2 => fsm_com_n_562, ZN => fsm_com_n_82);
  fsm_com_g21346 : ND2D1BWP7T port map(A1 => fsm_com_n_36, A2 => fsm_com_n_31, ZN => fsm_com_n_81);
  fsm_com_g21347 : CKND2D1BWP7T port map(A1 => yplayer(0), A2 => yplayer(1), ZN => fsm_com_n_79);
  fsm_com_g21348 : ND2D1BWP7T port map(A1 => level_abs(2), A2 => level_abs(0), ZN => fsm_com_n_78);
  fsm_com_g21349 : IND2D1BWP7T port map(A1 => xplayer(1), B1 => FE_PHN233_fsm_com_n_22, ZN => fsm_com_n_77);
  fsm_com_g21350 : ND2D1BWP7T port map(A1 => score_d(13), A2 => FE_PHN227_score_d_12, ZN => fsm_com_n_76);
  fsm_com_g21351 : ND2D1BWP7T port map(A1 => fsm_com_n_550, A2 => fsm_com_n_536, ZN => fsm_com_n_75);
  fsm_com_g21352 : NR2XD0BWP7T port map(A1 => energy_d(4), A2 => energy_d(5), ZN => fsm_com_n_74);
  fsm_com_g21353 : ND2D1BWP7T port map(A1 => fsm_com_n_549, A2 => fsm_com_n_571, ZN => fsm_com_n_73);
  fsm_com_g21354 : NR2D1BWP7T port map(A1 => fsm_com_n_538, A2 => FE_OFN0_reset, ZN => fsm_com_n_71);
  fsm_com_g21355 : NR2XD0BWP7T port map(A1 => fsm_com_n_555, A2 => fsm_com_n_561, ZN => fsm_com_n_70);
  fsm_com_g21356 : NR2XD0BWP7T port map(A1 => fsm_com_n_35, A2 => fsm_com_n_536, ZN => fsm_com_n_68);
  fsm_com_g21357 : NR2XD0BWP7T port map(A1 => fsm_com_n_560, A2 => fsm_com_n_563, ZN => fsm_com_n_66);
  fsm_com_g21358 : CKND1BWP7T port map(I => fsm_com_n_60, ZN => fsm_com_n_61);
  fsm_com_g21360 : INVD1BWP7T port map(I => fsm_com_n_52, ZN => fsm_com_n_53);
  fsm_com_g21361 : INVD0BWP7T port map(I => fsm_com_n_51, ZN => fsm_com_n_50);
  fsm_com_g21363 : INVD0BWP7T port map(I => fsm_com_n_44, ZN => fsm_com_n_43);
  fsm_com_g21364 : INVD0BWP7T port map(I => fsm_com_n_42, ZN => fsm_com_n_41);
  fsm_com_g21365 : NR2D1BWP7T port map(A1 => fsm_com_n_548, A2 => yplayer(0), ZN => fsm_com_n_40);
  fsm_com_g21366 : NR2D0BWP7T port map(A1 => fsm_com_n_572, A2 => map_data(18), ZN => fsm_com_n_39);
  fsm_com_g21367 : INR2XD0BWP7T port map(A1 => button_down, B1 => button_up, ZN => fsm_com_n_38);
  fsm_com_g21368 : OR2D0BWP7T port map(A1 => map_data(18), A2 => map_data(20), Z => fsm_com_n_63);
  fsm_com_g21369 : NR2XD0BWP7T port map(A1 => fsm_com_energy(0), A2 => fsm_com_energy(1), ZN => fsm_com_n_62);
  fsm_com_g21370 : NR2XD0BWP7T port map(A1 => map_data(38), A2 => map_data(36), ZN => fsm_com_n_60);
  fsm_com_g21371 : NR2XD0BWP7T port map(A1 => button_up, A2 => button_right, ZN => fsm_com_n_59);
  fsm_com_g21372 : NR2XD0BWP7T port map(A1 => fsm_com_n_548, A2 => fsm_com_n_547, ZN => fsm_com_n_58);
  fsm_com_g21373 : ND2D1BWP7T port map(A1 => level_d(1), A2 => level_d(0), ZN => fsm_com_n_57);
  fsm_com_g21374 : ND2D1BWP7T port map(A1 => level_d(5), A2 => level_d(4), ZN => fsm_com_n_56);
  fsm_com_g21375 : NR2D1BWP7T port map(A1 => fsm_com_n_29, A2 => fsm_com_n_571, ZN => fsm_com_n_55);
  fsm_com_g21376 : NR2XD0BWP7T port map(A1 => fsm_com_n_548, A2 => fsm_com_n_549, ZN => fsm_com_n_54);
  fsm_com_g21377 : NR2XD0BWP7T port map(A1 => level_abs(4), A2 => fsm_com_reached_high(1), ZN => fsm_com_n_52);
  fsm_com_g21378 : ND2D1BWP7T port map(A1 => xplayer(1), A2 => xplayer(0), ZN => fsm_com_n_51);
  fsm_com_g21379 : ND2D1BWP7T port map(A1 => score_d(9), A2 => FE_PHN249_score_d_8, ZN => fsm_com_n_49);
  fsm_com_g21380 : NR2XD0BWP7T port map(A1 => energy_d(8), A2 => energy_d(9), ZN => fsm_com_n_48);
  fsm_com_g21381 : NR2D1BWP7T port map(A1 => fsm_com_n_7, A2 => fsm_com_n_5, ZN => fsm_com_n_47);
  fsm_com_g21382 : NR2D1BWP7T port map(A1 => fsm_com_n_551, A2 => fsm_com_n_556, ZN => fsm_com_n_46);
  fsm_com_g21383 : CKND2D1BWP7T port map(A1 => fsm_com_n_547, A2 => fsm_com_n_565, ZN => fsm_com_n_44);
  fsm_com_g21384 : NR2D1BWP7T port map(A1 => fsm_com_n_33, A2 => fsm_com_n_565, ZN => fsm_com_n_42);
  fsm_com_g21450 : INVD1BWP7T port map(I => fsm_com_n_538, ZN => fsm_com_n_37);
  fsm_com_g21461 : INVD1BWP7T port map(I => fsm_com_n_557, ZN => fsm_com_n_36);
  fsm_com_g21462 : INVD1BWP7T port map(I => fsm_com_n_550, ZN => fsm_com_n_35);
  fsm_com_g21513 : INVD0BWP7T port map(I => fsm_com_n_547, ZN => fsm_com_n_33);
  fsm_com_g21530 : INVD0BWP7T port map(I => fsm_com_n_561, ZN => fsm_com_n_32);
  fsm_com_g21533 : INVD1BWP7T port map(I => fsm_com_n_555, ZN => fsm_com_n_31);
  fsm_com_g21534 : INVD1BWP7T port map(I => fsm_com_n_548, ZN => fsm_com_n_30);
  fsm_com_g21536 : INVD1BWP7T port map(I => fsm_com_n_549, ZN => fsm_com_n_29);
  fsm_com_energy_d_out_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => fsm_com_n_378, Q => FE_PHN247_energy_d_0, QN => fsm_com_n_5);
  fsm_com_energy_d_out_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => fsm_com_n_469, Q => FE_PHN246_energy_d_1, QN => fsm_com_n_7);
  fsm_com_energy_d_out_reg_2 : DFD1BWP7T port map(CP => CTS_20, D => fsm_com_n_479, Q => energy_d(2), QN => fsm_com_n_13);
  fsm_com_energy_d_out_reg_6 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN316_fsm_com_n_491, Q => energy_d(6), QN => fsm_com_n_18);
  fsm_com_energy_d_out_reg_10 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN502_fsm_com_n_489, Q => energy_d(10), QN => fsm_com_n_19);
  fsm_com_energy_reg_1 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_406, Q => fsm_com_energy(1), QN => fsm_com_n_4);
  fsm_com_energy_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => fsm_com_n_423, Q => fsm_com_energy(2), QN => fsm_com_n_15);
  fsm_com_energy_reg_4 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_409, Q => fsm_com_energy(4), QN => fsm_com_n_24);
  fsm_com_energy_reg_5 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN360_fsm_com_n_497, Q => fsm_com_energy(5), QN => fsm_com_n_26);
  fsm_com_energy_reg_6 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN355_fsm_com_n_482, Q => fsm_com_energy(6), QN => fsm_com_n_9);
  fsm_com_energy_reg_7 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_594, Q => fsm_com_energy(7), QN => fsm_com_n_23);
  fsm_com_level_reg_0 : DFD1BWP7T port map(CP => CTS_19, D => fsm_com_n_263, Q => FE_PHN243_level_abs_0, QN => fsm_com_n_16);
  fsm_com_level_reg_1 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN317_fsm_com_n_202, Q => level_abs(1), QN => fsm_com_n_21);
  fsm_com_level_reg_2 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_197, Q => level_abs(2), QN => fsm_com_n_25);
  fsm_com_level_reg_4 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN357_fsm_com_n_298, Q => level_abs(4), QN => fsm_com_n_14);
  fsm_com_score_d_out_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => fsm_com_n_428, Q => score_d(0), QN => fsm_com_n_28);
  fsm_com_score_d_out_reg_2 : DFD1BWP7T port map(CP => CTS_20, D => fsm_com_n_427, Q => score_d(2), QN => fsm_com_n_27);
  fsm_com_score_d_out_reg_3 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN262_fsm_com_n_434, Q => score_d(3), QN => fsm_com_n_17);
  fsm_com_x_pos_reg_0 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_331, Q => xplayer(0), QN => fsm_com_n_22);
  fsm_com_x_pos_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => fsm_com_n_369, Q => xplayer(2), QN => fsm_com_n_6);
  fsm_com_x_pos_reg_3 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_342, Q => xplayer(3), QN => FE_PHN365_fsm_com_n_20);
  fsm_com_y_pos_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => fsm_com_n_393, Q => yplayer(0), QN => fsm_com_n_11);
  fsm_com_y_pos_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => fsm_com_n_404, Q => yplayer(1), QN => fsm_com_n_8);
  fsm_com_y_pos_reg_2 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => fsm_com_n_396, Q => yplayer(2), QN => fsm_com_n_10);
  fsm_com_g2 : IND2D1BWP7T port map(A1 => fsm_com_n_402, B1 => fsm_com_n_152, ZN => fsm_com_n_3);
  fsm_com_g21585 : INR3D0BWP7T port map(A1 => fsm_com_n_284, B1 => fsm_com_n_415, B2 => fsm_com_n_166, ZN => fsm_com_n_2);
  fsm_com_g21586 : IND2D1BWP7T port map(A1 => fsm_com_n_171, B1 => fsm_com_n_132, ZN => fsm_com_n_1);
  fsm_com_g21587 : INR4D0BWP7T port map(A1 => fsm_com_n_59, B1 => button_down, B2 => button_left, B3 => button_mining, ZN => fsm_com_n_0);
  fsm_com_g21589 : ND3D0BWP7T port map(A1 => fsm_com_n_445, A2 => fsm_com_n_324, A3 => fsm_com_n_118, ZN => fsm_com_n_594);
  fsm_com_g21590 : INR2D1BWP7T port map(A1 => fsm_com_n_451, B1 => fsm_com_n_94, ZN => fsm_com_n_595);
  fsm_com_g21591 : IINR4D0BWP7T port map(A1 => fsm_com_n_375, A2 => fsm_com_n_299, B1 => fsm_com_n_66, B2 => fsm_com_n_543, ZN => fsm_com_n_596);
  fsm_com_g21592 : ND3D0BWP7T port map(A1 => fsm_com_n_386, A2 => fsm_com_n_320, A3 => fsm_com_n_116, ZN => fsm_com_n_597);
  fsm_com_g21593 : NR2D1BWP7T port map(A1 => fsm_com_n_391, A2 => fsm_com_n_310, ZN => fsm_com_n_598);
  fsm_com_g21594 : NR2D1BWP7T port map(A1 => fsm_com_n_309, A2 => fsm_com_n_47, ZN => fsm_com_n_599);
  fsm_com_g21595 : AN2D1BWP7T port map(A1 => fsm_com_n_244, A2 => fsm_com_n_211, Z => fsm_com_n_600);
  fsm_com_g21596 : ND2D1BWP7T port map(A1 => fsm_com_n_248, A2 => fsm_com_n_228, ZN => fsm_com_n_601);
  fsm_com_g21597 : IND2D1BWP7T port map(A1 => fsm_com_n_539, B1 => fsm_com_n_559, ZN => fsm_com_n_602);
  fsm_com_g21598 : IND2D1BWP7T port map(A1 => animation_done, B1 => fsm_com_n_546, ZN => fsm_com_n_603);
  fsm_com_g21599 : ND2D1BWP7T port map(A1 => fsm_com_n_567, A2 => fsm_com_n_548, ZN => fsm_com_n_604);
  fsm_com_score_d_out_reg_5 : DFD1BWP7T port map(CP => CTS_22, D => FE_PHN304_fsm_com_n_477, Q => score_d(5), QN => FE_PHN143_fsm_com_n_12);
  fsm_com_g21602 : AO21D0BWP7T port map(A1 => fsm_com_n_605, A2 => FE_PHN396_fsm_com_reached_high_0, B => fsm_com_n_322, Z => fsm_com_n_606);
  fsm_com_g3 : IND2D1BWP7T port map(A1 => fsm_com_n_286, B1 => fsm_com_n_214, ZN => fsm_com_n_605);
  vga_com_texture_module_g6969 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_vvis(5), A2 => vga_com_texture_module_n_663, B => vga_com_texture_module_n_664, ZN => vga_com_texture_module_n_703);
  vga_com_texture_module_g6971 : ND2D0BWP7T port map(A1 => vga_com_texture_module_vvis(5), A2 => vga_com_texture_module_n_663, ZN => vga_com_texture_module_n_664);
  vga_com_texture_module_g6972 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_9, A2 => vga_com_texture_module_n_662, B => vga_com_texture_module_n_663, Z => vga_com_texture_module_n_702);
  vga_com_texture_module_g6973 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_9, A2 => vga_com_texture_module_n_662, ZN => vga_com_texture_module_n_663);
  vga_com_texture_module_g6974 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_hvis(5), A2 => vga_com_texture_module_n_661, B => vga_com_texture_module_n_659, ZN => vga_com_texture_module_n_710);
  vga_com_texture_module_g6975 : MOAI22D0BWP7T port map(A1 => FE_PHN251_vga_com_texture_module_hvis_3, A2 => vga_com_texture_module_n_657, B1 => FE_PHN251_vga_com_texture_module_hvis_3, B2 => vga_com_texture_module_n_657, ZN => vga_com_texture_module_n_708);
  vga_com_texture_module_g6976 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_vvis(3), A2 => vga_com_texture_module_n_656, B1 => vga_com_texture_module_vvis(3), B2 => vga_com_texture_module_n_656, ZN => vga_com_texture_module_n_701);
  vga_com_texture_module_g6977 : INR2XD0BWP7T port map(A1 => vga_com_texture_module_n_656, B1 => vga_com_texture_module_vvis(3), ZN => vga_com_texture_module_n_662);
  vga_com_texture_module_g6978 : CKXOR2D1BWP7T port map(A1 => vga_com_texture_module_hvis(6), A2 => vga_com_texture_module_n_659, Z => vga_com_texture_module_n_711);
  vga_com_texture_module_g6979 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_hvis(4), A2 => vga_com_texture_module_n_658, B => vga_com_texture_module_n_660, ZN => vga_com_texture_module_n_709);
  vga_com_texture_module_g6980 : INVD0BWP7T port map(I => vga_com_texture_module_n_660, ZN => vga_com_texture_module_n_661);
  vga_com_texture_module_g6981 : CKND2D1BWP7T port map(A1 => vga_com_texture_module_hvis(4), A2 => vga_com_texture_module_n_658, ZN => vga_com_texture_module_n_660);
  vga_com_texture_module_g6982 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_670, B1 => vga_com_texture_module_n_658, ZN => vga_com_texture_module_n_659);
  vga_com_texture_module_g6983 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_vvis(2), A2 => vga_com_texture_module_n_654, B1 => vga_com_texture_module_vvis(2), B2 => vga_com_texture_module_n_654, ZN => vga_com_texture_module_n_700);
  vga_com_texture_module_g6984 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_hvis(2), A2 => vga_com_texture_module_n_655, B1 => vga_com_texture_module_hvis(2), B2 => vga_com_texture_module_n_655, ZN => vga_com_texture_module_n_707);
  vga_com_texture_module_g6985 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_675, A2 => vga_com_texture_module_n_655, ZN => vga_com_texture_module_n_658);
  vga_com_texture_module_g6986 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_655, B1 => vga_com_texture_module_hvis(2), ZN => vga_com_texture_module_n_657);
  vga_com_texture_module_g6987 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_654, B1 => vga_com_texture_module_vvis(2), ZN => vga_com_texture_module_n_656);
  vga_com_texture_module_g6988 : FA1D0BWP7T port map(A => vga_com_texture_module_n_652, B => vga_com_timer1(5), CI => vga_com_texture_module_n_650, CO => vga_com_texture_module_n_655, S => vga_com_texture_module_n_706);
  vga_com_texture_module_g6989 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_vvis(1), A2 => vga_com_texture_module_n_653, B1 => vga_com_texture_module_vvis(1), B2 => vga_com_texture_module_n_653, ZN => vga_com_texture_module_n_699);
  vga_com_texture_module_g6990 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_653, B1 => vga_com_texture_module_vvis(1), ZN => vga_com_texture_module_n_654);
  vga_com_texture_module_g6991 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_hvis(0), A2 => vga_com_texture_module_n_651, B => vga_com_texture_module_n_652, ZN => vga_com_texture_module_n_705);
  vga_com_texture_module_g6992 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_vvis(0), A2 => vga_com_texture_module_n_651, B => vga_com_texture_module_n_653, ZN => vga_com_texture_module_n_698);
  vga_com_texture_module_g6993 : CKND2D1BWP7T port map(A1 => vga_com_texture_module_vvis(4), A2 => vga_com_texture_module_vvis(5), ZN => vga_com_texture_module_n_671);
  vga_com_texture_module_g6994 : ND2D1BWP7T port map(A1 => vga_com_texture_module_hvis(4), A2 => vga_com_texture_module_hvis(5), ZN => vga_com_texture_module_n_670);
  vga_com_texture_module_g6995 : NR2XD0BWP7T port map(A1 => FE_PHN251_vga_com_texture_module_hvis_3, A2 => vga_com_texture_module_hvis(2), ZN => vga_com_texture_module_n_675);
  vga_com_texture_module_g6996 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_vvis(3), A2 => vga_com_texture_module_vvis(2), ZN => vga_com_texture_module_n_668);
  vga_com_texture_module_g6997 : ND2D1BWP7T port map(A1 => vga_com_texture_module_vvis(0), A2 => vga_com_texture_module_n_651, ZN => vga_com_texture_module_n_653);
  vga_com_texture_module_g6998 : ND2D1BWP7T port map(A1 => vga_com_texture_module_hvis(0), A2 => vga_com_texture_module_n_651, ZN => vga_com_texture_module_n_652);
  vga_com_texture_module_g16579 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_648, A2 => vga_com_texture_module_n_642, Z => vga_com_tile_address(1));
  vga_com_texture_module_g16580 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_648, A2 => vga_com_texture_module_n_636, Z => vga_com_tile_address(2));
  vga_com_texture_module_g16581 : OR3XD1BWP7T port map(A1 => vga_com_texture_module_n_269, A2 => vga_com_texture_module_n_645, A3 => vga_com_tile_address(3), Z => vga_com_texture_module_n_648);
  vga_com_texture_module_g16582 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_647, A2 => vga_com_texture_module_n_448, Z => vga_com_tile_address(3));
  vga_com_texture_module_g16583 : OAI31D0BWP7T port map(A1 => vga_com_texture_module_n_285, A2 => vga_com_texture_module_n_273, A3 => vga_com_texture_module_n_414, B => vga_com_texture_module_n_646, ZN => vga_com_texture_module_n_647);
  vga_com_texture_module_g16584 : AOI211D1BWP7T port map(A1 => vga_com_texture_module_n_449, A2 => vga_com_texture_module_frame_count(2), B => vga_com_texture_module_n_644, C => vga_com_texture_module_n_479, ZN => vga_com_texture_module_n_646);
  vga_com_texture_module_g16585 : IND4D0BWP7T port map(A1 => vga_com_tile_address(4), B1 => vga_com_texture_module_n_636, B2 => FE_OFN2_vga_com_tile_address_0, B3 => vga_com_texture_module_n_642, ZN => vga_com_texture_module_n_645);
  vga_com_texture_module_g16586 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_463, A2 => vga_com_texture_module_n_462, A3 => vga_com_texture_module_n_461, A4 => vga_com_texture_module_n_643, ZN => vga_com_texture_module_n_644);
  vga_com_texture_module_g16587 : AOI221D0BWP7T port map(A1 => vga_com_texture_module_n_424, A2 => energy_d(3), B1 => vga_com_texture_module_n_413, B2 => vga_com_texture_module_n_341, C => vga_com_texture_module_n_641, ZN => vga_com_texture_module_n_643);
  vga_com_texture_module_g16588 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_626, A2 => vga_com_texture_module_n_581, A3 => vga_com_texture_module_n_580, A4 => vga_com_texture_module_n_640, ZN => vga_com_texture_module_n_642);
  vga_com_texture_module_g16589 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_638, B1 => vga_com_texture_module_n_417, B2 => vga_com_texture_module_n_390, B3 => vga_com_texture_module_n_418, ZN => vga_com_texture_module_n_641);
  vga_com_texture_module_g16590 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_541, A2 => map_data(4), B => vga_com_texture_module_n_639, C => vga_com_texture_module_n_631, ZN => vga_com_texture_module_n_640);
  vga_com_texture_module_g16591 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_448, B1 => vga_com_texture_module_n_468, B2 => vga_com_texture_module_n_502, B3 => vga_com_texture_module_n_637, ZN => vga_com_texture_module_n_639);
  vga_com_texture_module_g16592 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_637, A2 => vga_com_texture_module_n_434, A3 => vga_com_texture_module_n_397, A4 => vga_com_texture_module_n_480, ZN => vga_com_texture_module_n_638);
  vga_com_texture_module_g16593 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_635, A2 => vga_com_texture_module_n_594, A3 => vga_com_texture_module_n_599, ZN => vga_com_texture_module_n_637);
  vga_com_texture_module_g16594 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_448, B1 => vga_com_texture_module_n_634, B2 => vga_com_texture_module_n_575, B3 => vga_com_texture_module_n_565, ZN => vga_com_texture_module_n_636);
  vga_com_texture_module_g16595 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_633, A2 => vga_com_texture_module_n_269, B1 => vga_com_texture_module_n_354, B2 => vga_com_texture_module_n_315, ZN => vga_com_texture_module_n_635);
  vga_com_texture_module_g16596 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_625, A2 => vga_com_texture_module_n_606, A3 => vga_com_texture_module_n_603, A4 => vga_com_texture_module_n_632, ZN => vga_com_tile_address(0));
  vga_com_texture_module_g16597 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_543, A2 => map_data(11), B => vga_com_texture_module_n_630, C => vga_com_texture_module_n_629, ZN => vga_com_texture_module_n_634);
  vga_com_texture_module_g16598 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_609, A2 => vga_com_texture_module_n_520, B => vga_com_texture_module_n_627, C => vga_com_texture_module_n_600, ZN => vga_com_texture_module_n_633);
  vga_com_texture_module_g16599 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_544, A2 => map_data(21), B => vga_com_texture_module_n_610, C => vga_com_texture_module_n_628, ZN => vga_com_texture_module_n_632);
  vga_com_texture_module_g16600 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_449, B1 => vga_com_texture_module_n_624, B2 => vga_com_texture_module_n_577, ZN => vga_com_texture_module_n_631);
  vga_com_texture_module_g16601 : OAI211D1BWP7T port map(A1 => vga_com_texture_module_n_340, A2 => vga_com_texture_module_n_390, B => vga_com_texture_module_n_623, C => vga_com_texture_module_n_601, ZN => vga_com_texture_module_n_630);
  vga_com_texture_module_g16602 : OR4D1BWP7T port map(A1 => vga_com_texture_module_n_484, A2 => vga_com_texture_module_n_481, A3 => vga_com_texture_module_n_619, A4 => vga_com_texture_module_n_612, Z => vga_com_texture_module_n_629);
  vga_com_texture_module_g16603 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_616, B1 => vga_com_texture_module_n_602, B2 => vga_com_texture_module_n_583, B3 => vga_com_texture_module_n_584, ZN => vga_com_texture_module_n_628);
  vga_com_texture_module_g16604 : OAI32D1BWP7T port map(A1 => vga_com_texture_module_n_333, A2 => vga_com_texture_module_n_324, A3 => vga_com_texture_module_n_345, B1 => vga_com_texture_module_n_344, B2 => vga_com_texture_module_n_620, ZN => vga_com_texture_module_n_627);
  vga_com_texture_module_g16605 : AOI221D0BWP7T port map(A1 => vga_com_texture_module_n_539, A2 => map_data(19), B1 => vga_com_texture_module_n_542, B2 => map_data(7), C => vga_com_texture_module_n_622, ZN => vga_com_texture_module_n_626);
  vga_com_texture_module_g16606 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_558, A2 => map_data(57), B => vga_com_texture_module_n_621, ZN => vga_com_texture_module_n_625);
  vga_com_texture_module_g16607 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_415, A2 => vga_com_texture_module_n_371, B => vga_com_texture_module_n_618, C => vga_com_texture_module_n_471, ZN => vga_com_texture_module_n_624);
  vga_com_texture_module_g16608 : AN4D1BWP7T port map(A1 => vga_com_texture_module_n_617, A2 => vga_com_texture_module_n_467, A3 => vga_com_texture_module_n_459, A4 => vga_com_texture_module_n_466, Z => vga_com_texture_module_n_623);
  vga_com_texture_module_g16609 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_559, A2 => map_data(67), B => vga_com_texture_module_n_615, Z => vga_com_texture_module_n_622);
  vga_com_texture_module_g16610 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_614, A2 => vga_com_texture_module_n_452, A3 => vga_com_texture_module_n_456, A4 => vga_com_texture_module_n_464, ZN => vga_com_texture_module_n_621);
  vga_com_texture_module_g16611 : AOI222D0BWP7T port map(A1 => vga_com_texture_module_n_609, A2 => vga_com_texture_module_n_570, B1 => vga_com_texture_module_n_571, B2 => vga_com_texture_module_n_513, C1 => vga_com_texture_module_n_535, C2 => vga_com_texture_module_n_515, ZN => vga_com_texture_module_n_620);
  vga_com_texture_module_g16612 : AO221D0BWP7T port map(A1 => vga_com_texture_module_n_540, A2 => map_data(17), B1 => vga_com_texture_module_n_541, B2 => map_data(5), C => vga_com_texture_module_n_611, Z => vga_com_texture_module_n_619);
  vga_com_texture_module_g16613 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_607, A2 => vga_com_texture_module_n_576, A3 => vga_com_texture_module_n_597, A4 => vga_com_texture_module_n_564, ZN => vga_com_texture_module_n_618);
  vga_com_texture_module_g16614 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_421, A2 => score_d(14), B => vga_com_texture_module_n_608, C => vga_com_texture_module_n_470, ZN => vga_com_texture_module_n_617);
  vga_com_texture_module_g16615 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_449, B1 => vga_com_texture_module_n_458, B2 => vga_com_texture_module_n_567, B3 => vga_com_texture_module_n_582, ZN => vga_com_texture_module_n_616);
  vga_com_texture_module_g16616 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_566, A2 => vga_com_texture_module_n_579, A3 => vga_com_texture_module_n_604, A4 => vga_com_texture_module_n_578, ZN => vga_com_texture_module_n_615);
  vga_com_texture_module_g16617 : OAI211D1BWP7T port map(A1 => vga_com_texture_module_n_325, A2 => vga_com_texture_module_n_426, B => vga_com_texture_module_n_438, C => vga_com_texture_module_n_613, ZN => vga_com_tile_address(4));
  vga_com_texture_module_g16618 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_393, A2 => level_d(0), B => vga_com_texture_module_n_605, ZN => vga_com_texture_module_n_614);
  vga_com_texture_module_g16619 : NR4D0BWP7T port map(A1 => vga_com_texture_module_n_474, A2 => vga_com_texture_module_n_472, A3 => vga_com_texture_module_n_441, A4 => vga_com_texture_module_n_596, ZN => vga_com_texture_module_n_613);
  vga_com_texture_module_g16620 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_598, A2 => vga_com_texture_module_n_569, A3 => vga_com_texture_module_n_591, A4 => vga_com_texture_module_n_593, ZN => vga_com_texture_module_n_612);
  vga_com_texture_module_g16621 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_588, A2 => vga_com_texture_module_n_590, A3 => vga_com_texture_module_n_589, A4 => vga_com_texture_module_n_595, ZN => vga_com_texture_module_n_611);
  vga_com_texture_module_g16622 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_587, A2 => vga_com_texture_module_n_568, A3 => vga_com_texture_module_n_585, A4 => vga_com_texture_module_n_586, ZN => vga_com_texture_module_n_610);
  vga_com_texture_module_g16623 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_599, B1 => vga_com_texture_module_n_435, B2 => vga_com_texture_module_n_395, B3 => vga_com_texture_module_n_465, ZN => vga_com_texture_module_n_608);
  vga_com_texture_module_g16624 : AOI221D0BWP7T port map(A1 => vga_com_texture_module_n_555, A2 => map_data(49), B1 => vga_com_texture_module_n_560, B2 => map_data(61), C => vga_com_texture_module_n_437, ZN => vga_com_texture_module_n_607);
  vga_com_texture_module_g16625 : AOI221D0BWP7T port map(A1 => vga_com_texture_module_n_563, A2 => map_data(39), B1 => vga_com_texture_module_n_545, B2 => FE_PHN507_map_data_24, C => vga_com_texture_module_n_574, ZN => vga_com_texture_module_n_606);
  vga_com_texture_module_g16626 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_573, A2 => vga_com_texture_module_n_482, A3 => vga_com_texture_module_n_487, A4 => vga_com_texture_module_n_439, ZN => vga_com_texture_module_n_605);
  vga_com_texture_module_g16627 : AN3D0BWP7T port map(A1 => vga_com_texture_module_n_571, A2 => vga_com_texture_module_n_530, A3 => vga_com_texture_module_n_537, Z => vga_com_texture_module_n_609);
  vga_com_texture_module_g16628 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_572, A2 => map_data(43), B1 => vga_com_texture_module_n_558, B2 => map_data(58), ZN => vga_com_texture_module_n_604);
  vga_com_texture_module_g16629 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_572, A2 => map_data(42), B1 => vga_com_texture_module_n_543, B2 => map_data(9), ZN => vga_com_texture_module_n_603);
  vga_com_texture_module_g16630 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_413, A2 => vga_com_texture_module_n_405, B => vga_com_texture_module_n_469, C => vga_com_texture_module_n_592, ZN => vga_com_texture_module_n_602);
  vga_com_texture_module_g16631 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_572, A2 => map_data(44), B1 => vga_com_texture_module_n_558, B2 => map_data(59), ZN => vga_com_texture_module_n_601);
  vga_com_texture_module_g16632 : AO22D0BWP7T port map(A1 => vga_com_texture_module_n_571, A2 => vga_com_texture_module_n_518, B1 => vga_com_texture_module_n_535, B2 => vga_com_texture_module_n_519, Z => vga_com_texture_module_n_600);
  vga_com_texture_module_g16633 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_556, A2 => map_data(56), B1 => vga_com_texture_module_n_559, B2 => map_data(68), ZN => vga_com_texture_module_n_598);
  vga_com_texture_module_g16634 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_561, A2 => map_data(46), B1 => vga_com_texture_module_n_420, B2 => vga_com_texture_module_n_402, ZN => vga_com_texture_module_n_597);
  vga_com_texture_module_g16635 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_551, A2 => vga_com_texture_module_n_381, A3 => vga_com_texture_module_n_488, A4 => vga_com_texture_module_n_486, ZN => vga_com_texture_module_n_596);
  vga_com_texture_module_g16636 : AOI32D1BWP7T port map(A1 => vga_com_texture_module_n_343, A2 => vga_com_texture_module_n_383, A3 => vga_com_texture_module_n_358, B1 => vga_com_texture_module_n_553, B2 => map_data(35), ZN => vga_com_texture_module_n_595);
  vga_com_texture_module_g16637 : OAI222D0BWP7T port map(A1 => vga_com_texture_module_n_547, A2 => vga_com_texture_module_n_389, B1 => vga_com_texture_module_n_355, B2 => vga_com_texture_module_n_365, C1 => vga_com_texture_module_n_345, C2 => vga_com_texture_module_n_302, ZN => vga_com_texture_module_n_594);
  vga_com_texture_module_g16638 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_554, A2 => map_data(53), B1 => vga_com_texture_module_n_539, B2 => map_data(20), ZN => vga_com_texture_module_n_593);
  vga_com_texture_module_g16639 : IOA21D1BWP7T port map(A1 => vga_com_texture_module_n_549, A2 => map_data(27), B => vga_com_texture_module_n_478, ZN => vga_com_texture_module_n_592);
  vga_com_texture_module_g16640 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_548, A2 => map_data(71), B1 => vga_com_texture_module_n_562, B2 => map_data(65), ZN => vga_com_texture_module_n_591);
  vga_com_texture_module_g16641 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_555, A2 => map_data(50), B1 => vga_com_texture_module_n_546, B2 => map_data(14), ZN => vga_com_texture_module_n_590);
  vga_com_texture_module_g16642 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_561, A2 => map_data(47), B1 => vga_com_texture_module_n_557, B2 => map_data(32), ZN => vga_com_texture_module_n_589);
  vga_com_texture_module_g16643 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_549, A2 => map_data(29), B1 => vga_com_texture_module_n_560, B2 => map_data(62), ZN => vga_com_texture_module_n_588);
  vga_com_texture_module_g16644 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_556, A2 => map_data(54), B1 => vga_com_texture_module_n_559, B2 => map_data(66), ZN => vga_com_texture_module_n_587);
  vga_com_texture_module_g16645 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_489, B1 => vga_com_texture_module_n_573, ZN => vga_com_texture_module_n_599);
  vga_com_texture_module_g16646 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_554, A2 => map_data(51), B1 => vga_com_texture_module_n_539, B2 => map_data(18), ZN => vga_com_texture_module_n_586);
  vga_com_texture_module_g16647 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_548, A2 => map_data(69), B1 => vga_com_texture_module_n_562, B2 => map_data(63), ZN => vga_com_texture_module_n_585);
  vga_com_texture_module_g16648 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_560, A2 => map_data(60), B1 => vga_com_texture_module_n_546, B2 => map_data(12), ZN => vga_com_texture_module_n_584);
  vga_com_texture_module_g16649 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_561, A2 => map_data(45), B1 => vga_com_texture_module_n_557, B2 => map_data(30), ZN => vga_com_texture_module_n_583);
  vga_com_texture_module_g16650 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_555, A2 => map_data(48), B1 => vga_com_texture_module_n_553, B2 => map_data(33), ZN => vga_com_texture_module_n_582);
  vga_com_texture_module_g16651 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_562, A2 => map_data(64), B1 => vga_com_texture_module_n_538, B2 => map_data(1), ZN => vga_com_texture_module_n_581);
  vga_com_texture_module_g16652 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_554, A2 => map_data(52), B1 => vga_com_texture_module_n_548, B2 => map_data(70), ZN => vga_com_texture_module_n_580);
  vga_com_texture_module_g16653 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_556, A2 => map_data(55), B1 => vga_com_texture_module_n_552, B2 => map_data(37), ZN => vga_com_texture_module_n_579);
  vga_com_texture_module_g16654 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_563, A2 => map_data(40), B1 => vga_com_texture_module_n_545, B2 => map_data(25), ZN => vga_com_texture_module_n_578);
  vga_com_texture_module_g16655 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_553, A2 => map_data(34), B1 => vga_com_texture_module_n_540, B2 => map_data(16), ZN => vga_com_texture_module_n_577);
  vga_com_texture_module_g16656 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_549, A2 => map_data(28), B1 => vga_com_texture_module_n_557, B2 => map_data(31), ZN => vga_com_texture_module_n_576);
  vga_com_texture_module_g16657 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_552, A2 => map_data(38), B1 => vga_com_texture_module_n_563, B2 => map_data(41), ZN => vga_com_texture_module_n_575);
  vga_com_texture_module_g16658 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_390, A2 => vga_com_texture_module_n_346, B1 => vga_com_texture_module_n_552, B2 => map_data(36), ZN => vga_com_texture_module_n_574);
  vga_com_texture_module_g16659 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_514, B1 => vga_com_texture_module_n_294, B2 => vga_com_texture_module_n_534, ZN => vga_com_texture_module_n_570);
  vga_com_texture_module_g16660 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_492, B1 => vga_com_texture_module_n_478, B2 => vga_com_texture_module_n_483, B3 => vga_com_texture_module_n_551, ZN => vga_com_tile_address(5));
  vga_com_texture_module_g16661 : AOI31D0BWP7T port map(A1 => vga_com_texture_module_n_678, A2 => vga_com_texture_module_n_356, A3 => vga_com_texture_module_n_401, B => vga_com_texture_module_n_550, ZN => vga_com_texture_module_n_573);
  vga_com_texture_module_g16662 : INR3D0BWP7T port map(A1 => vga_com_texture_module_n_519, B1 => vga_com_texture_module_n_269, B2 => vga_com_texture_module_n_535, ZN => vga_com_texture_module_n_572);
  vga_com_texture_module_g16663 : AN3D1BWP7T port map(A1 => vga_com_texture_module_n_532, A2 => vga_com_texture_module_n_536, A3 => vga_com_texture_module_n_535, Z => vga_com_texture_module_n_571);
  vga_com_texture_module_g16664 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_538, A2 => map_data(2), B1 => vga_com_texture_module_n_542, B2 => map_data(8), ZN => vga_com_texture_module_n_569);
  vga_com_texture_module_g16665 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_538, A2 => map_data(0), B1 => vga_com_texture_module_n_542, B2 => map_data(6), ZN => vga_com_texture_module_n_568);
  vga_com_texture_module_g16666 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_540, A2 => map_data(15), B1 => vga_com_texture_module_n_541, B2 => map_data(3), ZN => vga_com_texture_module_n_567);
  vga_com_texture_module_g16667 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_544, A2 => map_data(22), B1 => vga_com_texture_module_n_543, B2 => map_data(10), ZN => vga_com_texture_module_n_566);
  vga_com_texture_module_g16668 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_544, A2 => map_data(23), B1 => vga_com_texture_module_n_545, B2 => FE_PHN501_map_data_26, ZN => vga_com_texture_module_n_565);
  vga_com_texture_module_g16669 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_546, A2 => map_data(13), B1 => vga_com_texture_module_n_451, B2 => vga_com_texture_module_n_260, ZN => vga_com_texture_module_n_564);
  vga_com_texture_module_g16670 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_525, B1 => vga_com_texture_module_n_535, ZN => vga_com_texture_module_n_563);
  vga_com_texture_module_g16671 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_521, A2 => vga_com_texture_module_n_537, ZN => vga_com_texture_module_n_562);
  vga_com_texture_module_g16672 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_523, A2 => vga_com_texture_module_n_536, ZN => vga_com_texture_module_n_561);
  vga_com_texture_module_g16673 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_522, A2 => vga_com_texture_module_n_537, ZN => vga_com_texture_module_n_560);
  vga_com_texture_module_g16674 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_526, A2 => vga_com_texture_module_n_537, ZN => vga_com_texture_module_n_559);
  vga_com_texture_module_g16675 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_525, B1 => vga_com_texture_module_n_536, ZN => vga_com_texture_module_n_558);
  vga_com_texture_module_g16676 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_523, A2 => vga_com_texture_module_n_535, ZN => vga_com_texture_module_n_557);
  vga_com_texture_module_g16677 : NR2D0BWP7T port map(A1 => vga_com_texture_module_n_526, A2 => vga_com_texture_module_n_536, ZN => vga_com_texture_module_n_556);
  vga_com_texture_module_g16678 : INVD0BWP7T port map(I => vga_com_texture_module_n_550, ZN => vga_com_texture_module_n_551);
  vga_com_texture_module_g16679 : OR4XD1BWP7T port map(A1 => vga_com_texture_module_n_518, A2 => vga_com_texture_module_n_519, A3 => vga_com_texture_module_n_520, A4 => vga_com_texture_module_n_527, Z => vga_com_texture_module_n_547);
  vga_com_texture_module_g16680 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_522, A2 => vga_com_texture_module_n_536, ZN => vga_com_texture_module_n_555);
  vga_com_texture_module_g16681 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_521, A2 => vga_com_texture_module_n_536, ZN => vga_com_texture_module_n_554);
  vga_com_texture_module_g16682 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_522, A2 => vga_com_texture_module_n_535, ZN => vga_com_texture_module_n_553);
  vga_com_texture_module_g16683 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_526, A2 => vga_com_texture_module_n_535, ZN => vga_com_texture_module_n_552);
  vga_com_texture_module_g16684 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_521, A2 => vga_com_texture_module_n_535, ZN => vga_com_texture_module_n_550);
  vga_com_texture_module_g16685 : INR3D0BWP7T port map(A1 => vga_com_texture_module_n_515, B1 => vga_com_texture_module_n_389, B2 => vga_com_texture_module_n_535, ZN => vga_com_texture_module_n_549);
  vga_com_texture_module_g16686 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_521, A2 => vga_com_texture_module_n_531, A3 => vga_com_texture_module_n_376, ZN => vga_com_texture_module_n_548);
  vga_com_texture_module_g16687 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_523, A2 => vga_com_texture_module_n_532, ZN => vga_com_texture_module_n_546);
  vga_com_texture_module_g16688 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_525, B1 => vga_com_texture_module_n_532, ZN => vga_com_texture_module_n_545);
  vga_com_texture_module_g16689 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_526, A2 => vga_com_texture_module_n_532, ZN => vga_com_texture_module_n_544);
  vga_com_texture_module_g16690 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_526, A2 => vga_com_texture_module_n_530, ZN => vga_com_texture_module_n_543);
  vga_com_texture_module_g16691 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_521, A2 => vga_com_texture_module_n_530, ZN => vga_com_texture_module_n_542);
  vga_com_texture_module_g16692 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_522, A2 => vga_com_texture_module_n_530, ZN => vga_com_texture_module_n_541);
  vga_com_texture_module_g16693 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_529, A2 => vga_com_texture_module_n_375, B1 => vga_com_texture_module_n_524, B2 => vga_com_texture_module_n_376, ZN => vga_com_texture_module_n_534);
  vga_com_texture_module_g16694 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_522, A2 => vga_com_texture_module_n_532, ZN => vga_com_texture_module_n_540);
  vga_com_texture_module_g16695 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_521, A2 => vga_com_texture_module_n_532, ZN => vga_com_texture_module_n_539);
  vga_com_texture_module_g16696 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_521, A2 => vga_com_texture_module_n_528, A3 => vga_com_texture_module_n_375, ZN => vga_com_texture_module_n_538);
  vga_com_texture_module_g16697 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_376, B1 => vga_com_texture_module_n_533, ZN => vga_com_texture_module_n_537);
  vga_com_texture_module_g16698 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_531, B1 => vga_com_texture_module_n_376, ZN => vga_com_texture_module_n_536);
  vga_com_texture_module_g16699 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_533, A2 => vga_com_texture_module_n_376, ZN => vga_com_texture_module_n_535);
  vga_com_texture_module_g16700 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_529, A2 => vga_com_texture_module_n_294, ZN => vga_com_texture_module_n_533);
  vga_com_texture_module_g16701 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_528, A2 => vga_com_texture_module_n_376, Z => vga_com_texture_module_n_532);
  vga_com_texture_module_g16702 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_529, B1 => vga_com_texture_module_n_294, ZN => vga_com_texture_module_n_531);
  vga_com_texture_module_g16703 : OR3D1BWP7T port map(A1 => vga_com_texture_module_n_294, A2 => vga_com_texture_module_n_376, A3 => vga_com_texture_module_n_524, Z => vga_com_texture_module_n_530);
  vga_com_texture_module_g16704 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_504, A2 => vga_com_texture_module_n_512, A3 => vga_com_texture_module_n_498, ZN => vga_com_texture_module_n_529);
  vga_com_texture_module_g16705 : OR4XD1BWP7T port map(A1 => vga_com_texture_module_n_514, A2 => vga_com_texture_module_n_517, A3 => vga_com_texture_module_n_513, A4 => vga_com_texture_module_n_515, Z => vga_com_texture_module_n_527);
  vga_com_texture_module_g16706 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_524, B1 => vga_com_texture_module_n_294, ZN => vga_com_texture_module_n_528);
  vga_com_texture_module_g16707 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_520, A2 => vga_com_texture_module_n_268, ZN => vga_com_texture_module_n_526);
  vga_com_texture_module_g16708 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_518, A2 => vga_com_texture_module_n_268, Z => vga_com_texture_module_n_525);
  vga_com_texture_module_g16709 : OR3D1BWP7T port map(A1 => vga_com_texture_module_n_498, A2 => vga_com_texture_module_n_508, A3 => vga_com_texture_module_n_504, Z => vga_com_texture_module_n_524);
  vga_com_texture_module_g16710 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_389, B1 => vga_com_texture_module_n_513, ZN => vga_com_texture_module_n_523);
  vga_com_texture_module_g16711 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_389, B1 => vga_com_texture_module_n_514, ZN => vga_com_texture_module_n_522);
  vga_com_texture_module_g16712 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_389, B1 => vga_com_texture_module_n_517, ZN => vga_com_texture_module_n_521);
  vga_com_texture_module_g16713 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_516, A2 => vga_com_texture_module_n_377, ZN => vga_com_texture_module_n_520);
  vga_com_texture_module_g16714 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_516, A2 => vga_com_texture_module_n_378, ZN => vga_com_texture_module_n_519);
  vga_com_texture_module_g16715 : AN3D1BWP7T port map(A1 => vga_com_texture_module_n_510, A2 => vga_com_texture_module_n_378, A3 => vga_com_texture_module_n_295, Z => vga_com_texture_module_n_518);
  vga_com_texture_module_g16716 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_511, A2 => vga_com_texture_module_n_378, ZN => vga_com_texture_module_n_517);
  vga_com_texture_module_g16717 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_295, B1 => vga_com_texture_module_n_510, ZN => vga_com_texture_module_n_516);
  vga_com_texture_module_g16718 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_509, A2 => vga_com_texture_module_n_377, ZN => vga_com_texture_module_n_515);
  vga_com_texture_module_g16719 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_503, A2 => vga_com_texture_module_yposition(4), B => vga_com_texture_module_n_507, ZN => vga_com_texture_module_n_512);
  vga_com_texture_module_g16720 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_509, A2 => vga_com_texture_module_n_378, ZN => vga_com_texture_module_n_514);
  vga_com_texture_module_g16721 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_511, A2 => vga_com_texture_module_n_377, ZN => vga_com_texture_module_n_513);
  vga_com_texture_module_g16722 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_506, A2 => vga_com_texture_module_n_295, ZN => vga_com_texture_module_n_511);
  vga_com_texture_module_g16723 : NR4D0BWP7T port map(A1 => vga_com_texture_module_n_505, A2 => vga_com_texture_module_n_496, A3 => vga_com_texture_module_n_267, A4 => vga_com_texture_module_xposition(4), ZN => vga_com_texture_module_n_510);
  vga_com_texture_module_g16724 : INVD0BWP7T port map(I => vga_com_texture_module_n_507, ZN => vga_com_texture_module_n_508);
  vga_com_texture_module_g16725 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_295, B1 => vga_com_texture_module_n_506, ZN => vga_com_texture_module_n_509);
  vga_com_texture_module_g16726 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_503, A2 => vga_com_texture_module_yposition(4), ZN => vga_com_texture_module_n_507);
  vga_com_texture_module_g16727 : AN3D1BWP7T port map(A1 => vga_com_texture_module_n_505, A2 => vga_com_texture_module_n_496, A3 => vga_com_texture_module_n_282, Z => vga_com_texture_module_n_506);
  vga_com_texture_module_g16728 : AO211D0BWP7T port map(A1 => vga_com_texture_module_n_447, A2 => vga_com_texture_module_n_446, B => vga_com_dim(2), C => vga_com_texture_module_n_494, Z => vga_com_dim(1));
  vga_com_texture_module_g16729 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_500, A2 => vga_com_texture_module_xposition(3), B1 => vga_com_texture_module_n_500, B2 => vga_com_texture_module_xposition(3), ZN => vga_com_texture_module_n_505);
  vga_com_texture_module_g16730 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_501, A2 => yplayer(3), B1 => vga_com_texture_module_n_501, B2 => yplayer(3), ZN => vga_com_texture_module_n_504);
  vga_com_texture_module_g16731 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_499, A2 => vga_com_texture_module_n_491, B => vga_com_texture_module_n_485, ZN => vga_com_dim(2));
  vga_com_texture_module_g16732 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_457, A2 => vga_com_texture_module_n_346, B => vga_com_texture_module_n_493, C => vga_com_texture_module_n_453, ZN => vga_com_texture_module_n_502);
  vga_com_texture_module_g16733 : MAOI222D1BWP7T port map(A => vga_com_texture_module_n_497, B => vga_com_texture_module_n_25, C => yplayer(3), ZN => vga_com_texture_module_n_503);
  vga_com_texture_module_g16734 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_497, A2 => vga_com_texture_module_n_25, B1 => vga_com_texture_module_n_497, B2 => vga_com_texture_module_n_25, ZN => vga_com_texture_module_n_501);
  vga_com_texture_module_g16735 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_495, A2 => xplayer(3), B1 => vga_com_texture_module_n_495, B2 => xplayer(3), ZN => vga_com_texture_module_n_500);
  vga_com_texture_module_g16736 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_447, A2 => vga_com_texture_module_n_490, B => vga_com_texture_module_n_429, ZN => vga_com_texture_module_n_499);
  vga_com_texture_module_g16737 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_494, B1 => vga_com_texture_module_n_485, ZN => vga_com_dim(3));
  vga_com_texture_module_g16738 : FA1D0BWP7T port map(A => vga_com_texture_module_n_7, B => yplayer(2), CI => vga_com_texture_module_n_370, CO => vga_com_texture_module_n_497, S => vga_com_texture_module_n_498);
  vga_com_texture_module_g16739 : FA1D0BWP7T port map(A => vga_com_texture_module_n_259, B => xplayer(2), CI => vga_com_texture_module_n_369, CO => vga_com_texture_module_n_495, S => vga_com_texture_module_n_496);
  vga_com_texture_module_g16740 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_491, B1 => vga_com_texture_module_n_389, ZN => vga_com_texture_module_n_494);
  vga_com_texture_module_g16741 : ND4D0BWP7T port map(A1 => vga_com_texture_module_n_455, A2 => vga_com_texture_module_n_476, A3 => vga_com_texture_module_n_460, A4 => vga_com_texture_module_n_477, ZN => vga_com_texture_module_n_493);
  vga_com_texture_module_g16742 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_302, A2 => vga_com_texture_module_n_473, B1 => vga_com_texture_module_n_342, B2 => vga_com_texture_module_n_358, ZN => vga_com_texture_module_n_492);
  vga_com_texture_module_g16743 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_276, A2 => vga_com_texture_module_n_475, ZN => vga_com_texture_module_n_490);
  vga_com_texture_module_g16744 : AOI31D0BWP7T port map(A1 => vga_com_texture_module_n_409, A2 => vga_com_texture_module_n_351, A3 => vga_com_texture_module_n_319, B => vga_com_texture_module_n_302, ZN => vga_com_texture_module_n_489);
  vga_com_texture_module_g16745 : NR4D0BWP7T port map(A1 => vga_com_texture_module_n_403, A2 => vga_com_texture_module_n_411, A3 => vga_com_texture_module_n_443, A4 => vga_com_texture_module_n_440, ZN => vga_com_texture_module_n_488);
  vga_com_texture_module_g16746 : AOI221D0BWP7T port map(A1 => vga_com_texture_module_n_424, A2 => energy_d(0), B1 => vga_com_texture_module_n_423, B2 => energy_d(4), C => vga_com_texture_module_n_433, ZN => vga_com_texture_module_n_487);
  vga_com_texture_module_g16747 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_348, A2 => vga_com_texture_module_n_313, B => vga_com_texture_module_n_479, ZN => vga_com_texture_module_n_486);
  vga_com_texture_module_g16748 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_262, A2 => vga_com_texture_module_n_410, B => vga_com_texture_module_n_287, C => vga_com_texture_module_n_368, ZN => vga_com_texture_module_n_491);
  vga_com_texture_module_g16749 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_419, A2 => vga_com_texture_module_n_683, B1 => vga_com_texture_module_n_450, B2 => vga_com_texture_module_n_712, ZN => vga_com_texture_module_n_484);
  vga_com_texture_module_g16750 : AO211D0BWP7T port map(A1 => vga_com_texture_module_n_430, A2 => vga_com_texture_module_n_404, B => vga_com_texture_module_n_429, C => vga_com_texture_module_n_447, Z => vga_com_dim(0));
  vga_com_texture_module_g16751 : AOI32D1BWP7T port map(A1 => vga_com_texture_module_n_420, A2 => vga_com_texture_module_n_272, A3 => vga_com_texture_module_frame_count(3), B1 => vga_com_texture_module_n_413, B2 => vga_com_texture_module_n_366, ZN => vga_com_texture_module_n_483);
  vga_com_texture_module_g16752 : AOI222D0BWP7T port map(A1 => vga_com_texture_module_n_347, A2 => vga_com_texture_module_n_388, B1 => vga_com_texture_module_n_406, B2 => vga_com_texture_module_n_289, C1 => vga_com_texture_module_n_394, C2 => level_d(4), ZN => vga_com_texture_module_n_482);
  vga_com_texture_module_g16753 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_445, A2 => vga_com_texture_module_n_312, B1 => vga_com_texture_module_n_412, B2 => vga_com_texture_module_n_373, ZN => vga_com_texture_module_n_481);
  vga_com_texture_module_g16754 : AOI31D0BWP7T port map(A1 => vga_com_texture_module_n_392, A2 => vga_com_texture_module_n_356, A3 => vga_com_texture_module_n_329, B => vga_com_texture_module_n_454, ZN => vga_com_texture_module_n_480);
  vga_com_texture_module_g16755 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_429, A2 => vga_com_texture_module_n_444, B1 => vga_com_texture_module_n_287, B2 => vga_com_texture_module_n_431, ZN => vga_com_texture_module_n_485);
  vga_com_texture_module_g16756 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_423, A2 => energy_d(5), B1 => vga_com_texture_module_n_382, B2 => energy_d(9), ZN => vga_com_texture_module_n_477);
  vga_com_texture_module_g16757 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_428, A2 => score_d(9), B1 => vga_com_texture_module_n_421, B2 => score_d(13), ZN => vga_com_texture_module_n_476);
  vga_com_texture_module_g16758 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_407, A2 => vga_com_texture_module_n_691, B => vga_com_texture_module_n_693, ZN => vga_com_texture_module_n_475);
  vga_com_texture_module_g16759 : OAI31D0BWP7T port map(A1 => vga_com_texture_module_n_352, A2 => vga_com_texture_module_n_400, A3 => vga_com_texture_module_n_418, B => vga_com_texture_module_n_442, ZN => vga_com_texture_module_n_474);
  vga_com_texture_module_g16760 : AOI31D0BWP7T port map(A1 => vga_com_texture_module_n_345, A2 => vga_com_texture_module_n_349, A3 => vga_com_texture_module_n_316, B => vga_com_texture_module_n_436, ZN => vga_com_texture_module_n_473);
  vga_com_texture_module_g16761 : OA21D0BWP7T port map(A1 => vga_com_texture_module_n_347, A2 => vga_com_texture_module_n_432, B => vga_com_texture_module_n_355, Z => vga_com_texture_module_n_472);
  vga_com_texture_module_g16762 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_412, A2 => vga_com_texture_module_n_372, B1 => vga_com_texture_module_n_426, B2 => vga_com_texture_module_n_374, ZN => vga_com_texture_module_n_471);
  vga_com_texture_module_g16763 : AOI211D0BWP7T port map(A1 => vga_com_texture_module_n_356, A2 => vga_com_texture_module_n_352, B => vga_com_texture_module_n_417, C => vga_com_texture_module_n_357, ZN => vga_com_texture_module_n_470);
  vga_com_texture_module_g16764 : AOI31D0BWP7T port map(A1 => vga_com_texture_module_n_385, A2 => vga_com_texture_module_n_367, A3 => vga_com_texture_module_n_346, B => vga_com_texture_module_n_342, ZN => vga_com_texture_module_n_469);
  vga_com_texture_module_g16765 : AOI32D1BWP7T port map(A1 => vga_com_texture_module_n_392, A2 => vga_com_texture_module_n_386, A3 => vga_com_texture_module_n_360, B1 => vga_com_texture_module_n_393, B2 => level_d(1), ZN => vga_com_texture_module_n_468);
  vga_com_texture_module_g16766 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_428, A2 => score_d(10), B1 => vga_com_texture_module_n_422, B2 => score_d(6), ZN => vga_com_texture_module_n_467);
  vga_com_texture_module_g16767 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_424, A2 => energy_d(2), B1 => vga_com_texture_module_n_423, B2 => energy_d(6), ZN => vga_com_texture_module_n_466);
  vga_com_texture_module_g16768 : INR2D0BWP7T port map(A1 => vga_com_texture_module_n_285, B1 => vga_com_texture_module_n_450, ZN => vga_com_texture_module_n_479);
  vga_com_texture_module_g16769 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_676, B1 => vga_com_texture_module_n_451, ZN => vga_com_texture_module_n_478);
  vga_com_texture_module_g16770 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_392, A2 => vga_com_texture_module_n_323, B1 => vga_com_texture_module_n_418, B2 => vga_com_texture_module_n_317, ZN => vga_com_texture_module_n_465);
  vga_com_texture_module_g16771 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_427, A2 => score_d(0), B1 => vga_com_texture_module_n_382, B2 => energy_d(8), ZN => vga_com_texture_module_n_464);
  vga_com_texture_module_g16772 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_428, A2 => score_d(11), B1 => vga_com_texture_module_n_421, B2 => score_d(15), ZN => vga_com_texture_module_n_463);
  vga_com_texture_module_g16773 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_427, A2 => score_d(3), B1 => vga_com_texture_module_n_422, B2 => score_d(7), ZN => vga_com_texture_module_n_462);
  vga_com_texture_module_g16774 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_423, A2 => energy_d(7), B1 => vga_com_texture_module_n_382, B2 => energy_d(11), ZN => vga_com_texture_module_n_461);
  vga_com_texture_module_g16775 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_427, A2 => score_d(1), B1 => vga_com_texture_module_n_422, B2 => score_d(5), ZN => vga_com_texture_module_n_460);
  vga_com_texture_module_g16776 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_427, A2 => score_d(2), B1 => vga_com_texture_module_n_382, B2 => energy_d(10), ZN => vga_com_texture_module_n_459);
  vga_com_texture_module_g16777 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_425, A2 => vga_com_texture_module_n_325, B1 => vga_com_texture_module_n_415, B2 => vga_com_texture_module_n_339, ZN => vga_com_texture_module_n_458);
  vga_com_texture_module_g16778 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_417, A2 => vga_com_texture_module_n_318, B1 => vga_com_texture_module_n_390, B2 => vga_com_texture_module_n_322, ZN => vga_com_texture_module_n_457);
  vga_com_texture_module_g16779 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_421, A2 => score_d(12), B1 => vga_com_texture_module_n_418, B2 => vga_com_texture_module_n_321, ZN => vga_com_texture_module_n_456);
  vga_com_texture_module_g16780 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_424, A2 => FE_PHN403_energy_d_1, B1 => vga_com_texture_module_n_395, B2 => vga_com_texture_module_n_355, ZN => vga_com_texture_module_n_455);
  vga_com_texture_module_g16781 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_387, A2 => vga_com_texture_module_n_357, B1 => vga_com_texture_module_n_426, B2 => vga_com_texture_module_n_311, ZN => vga_com_texture_module_n_454);
  vga_com_texture_module_g16782 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_418, A2 => vga_com_texture_module_n_318, B1 => vga_com_texture_module_n_394, B2 => level_d(5), ZN => vga_com_texture_module_n_453);
  vga_com_texture_module_g16783 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_428, A2 => FE_PHN249_score_d_8, B1 => vga_com_texture_module_n_422, B2 => FE_PHN244_score_d_4, ZN => vga_com_texture_module_n_452);
  vga_com_texture_module_g16784 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_692, B1 => vga_com_texture_module_n_326, B2 => vga_com_texture_module_n_277, B3 => vga_com_texture_module_n_368, ZN => vga_com_texture_module_n_446);
  vga_com_texture_module_g16785 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_415, A2 => vga_com_texture_module_n_396, ZN => vga_com_texture_module_n_445);
  vga_com_texture_module_g16786 : AO211D0BWP7T port map(A1 => vga_com_texture_module_n_275, A2 => vga_com_texture_module_n_337, B => vga_com_texture_module_n_697, C => vga_com_texture_module_n_694, Z => vga_com_texture_module_n_444);
  vga_com_texture_module_g16787 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_399, A2 => vga_com_texture_module_n_398, B => vga_com_texture_module_n_269, ZN => vga_com_texture_module_n_443);
  vga_com_texture_module_g16788 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_356, A2 => vga_com_texture_module_n_358, B => vga_com_texture_module_n_417, Z => vga_com_texture_module_n_442);
  vga_com_texture_module_g16789 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_419, A2 => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_451);
  vga_com_texture_module_g16790 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_413, A2 => vga_com_texture_module_n_273, ZN => vga_com_texture_module_n_450);
  vga_com_texture_module_g16791 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_414, A2 => vga_com_texture_module_n_263, ZN => vga_com_texture_module_n_449);
  vga_com_texture_module_g16792 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_432, A2 => vga_com_texture_module_n_356, Z => vga_com_texture_module_n_448);
  vga_com_texture_module_g16793 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_694, B1 => vga_com_texture_module_n_431, ZN => vga_com_texture_module_n_447);
  vga_com_texture_module_g16794 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_385, A2 => vga_com_texture_module_n_360, B => vga_com_texture_module_n_342, ZN => vga_com_texture_module_n_441);
  vga_com_texture_module_g16795 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_362, A2 => vga_com_texture_module_frame_count(3), B => vga_com_texture_module_n_414, ZN => vga_com_texture_module_n_440);
  vga_com_texture_module_g16796 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_400, A2 => vga_com_texture_module_n_357, B => vga_com_texture_module_n_416, ZN => vga_com_texture_module_n_439);
  vga_com_texture_module_g16797 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_387, A2 => vga_com_texture_module_n_390, B => vga_com_texture_module_n_346, Z => vga_com_texture_module_n_438);
  vga_com_texture_module_g16798 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_383, A2 => vga_com_texture_module_n_346, B => vga_com_texture_module_n_342, ZN => vga_com_texture_module_n_437);
  vga_com_texture_module_g16799 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_316, A2 => vga_com_texture_module_n_332, B => vga_com_texture_module_n_408, ZN => vga_com_texture_module_n_436);
  vga_com_texture_module_g16800 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_393, A2 => level_d(2), B1 => vga_com_texture_module_n_394, B2 => level_d(6), ZN => vga_com_texture_module_n_435);
  vga_com_texture_module_g16801 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_393, A2 => level_d(3), B1 => vga_com_texture_module_n_394, B2 => level_d(7), ZN => vga_com_texture_module_n_434);
  vga_com_texture_module_g16802 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_283, A2 => vga_com_texture_module_n_681, B1 => vga_com_texture_module_n_28, B2 => vga_com_texture_module_n_683, ZN => animation_done);
  vga_com_texture_module_g16803 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_391, A2 => vga_com_texture_module_n_386, B1 => vga_com_texture_module_n_302, B2 => vga_com_texture_module_n_351, ZN => vga_com_texture_module_n_433);
  vga_com_texture_module_g16804 : INVD0BWP7T port map(I => vga_com_texture_module_n_431, ZN => vga_com_texture_module_n_430);
  vga_com_texture_module_g16805 : INVD0BWP7T port map(I => vga_com_texture_module_n_426, ZN => vga_com_texture_module_n_425);
  vga_com_texture_module_g16806 : CKND1BWP7T port map(I => vga_com_texture_module_n_420, ZN => vga_com_texture_module_n_419);
  vga_com_texture_module_g16807 : AN2D0BWP7T port map(A1 => vga_com_texture_module_n_289, A2 => vga_com_texture_module_n_401, Z => vga_com_texture_module_n_432);
  vga_com_texture_module_g16808 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_389, B1 => vga_com_texture_module_n_695, ZN => vga_com_texture_module_n_431);
  vga_com_texture_module_g16809 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_287, A2 => vga_com_texture_module_n_389, ZN => vga_com_texture_module_n_429);
  vga_com_texture_module_g16810 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_380, A2 => vga_com_texture_module_n_329, ZN => vga_com_texture_module_n_428);
  vga_com_texture_module_g16811 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_379, A2 => vga_com_texture_module_n_363, Z => vga_com_texture_module_n_427);
  vga_com_texture_module_g16812 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_396, A2 => vga_com_texture_module_n_355, ZN => vga_com_texture_module_n_426);
  vga_com_texture_module_g16813 : NR2D0BWP7T port map(A1 => vga_com_texture_module_n_269, A2 => vga_com_texture_module_n_399, ZN => vga_com_texture_module_n_424);
  vga_com_texture_module_g16814 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_269, A2 => vga_com_texture_module_n_398, ZN => vga_com_texture_module_n_423);
  vga_com_texture_module_g16815 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_380, A2 => vga_com_texture_module_n_359, ZN => vga_com_texture_module_n_422);
  vga_com_texture_module_g16816 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_380, A2 => vga_com_texture_module_n_330, ZN => vga_com_texture_module_n_421);
  vga_com_texture_module_g16817 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_397, A2 => vga_com_texture_module_n_356, ZN => vga_com_texture_module_n_420);
  vga_com_texture_module_g16818 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_379, A2 => vga_com_texture_module_n_384, ZN => vga_com_texture_module_n_418);
  vga_com_texture_module_g16819 : INVD0BWP7T port map(I => vga_com_texture_module_n_416, ZN => vga_com_texture_module_n_417);
  vga_com_texture_module_g16820 : INVD0BWP7T port map(I => vga_com_texture_module_n_415, ZN => vga_com_texture_module_n_414);
  vga_com_texture_module_g16821 : INVD0BWP7T port map(I => vga_com_texture_module_n_413, ZN => vga_com_texture_module_n_412);
  vga_com_texture_module_g16822 : NR2D0BWP7T port map(A1 => vga_com_texture_module_n_380, A2 => vga_com_texture_module_n_384, ZN => vga_com_texture_module_n_411);
  vga_com_texture_module_g16823 : OAI31D0BWP7T port map(A1 => vga_com_texture_module_n_334, A2 => vga_com_texture_module_n_689, A3 => vga_com_texture_module_n_690, B => vga_com_texture_module_n_692, ZN => vga_com_texture_module_n_410);
  vga_com_texture_module_g16824 : AOI222D0BWP7T port map(A1 => vga_com_texture_module_n_335, A2 => vga_com_texture_module_n_265, B1 => vga_com_texture_module_n_310, B2 => vga_com_texture_module_n_270, C1 => vga_com_texture_module_n_296, C2 => vga_com_texture_module_xposition(0), ZN => vga_com_texture_module_n_409);
  vga_com_texture_module_g16825 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_349, B1 => vga_com_texture_module_n_329, B2 => vga_com_texture_module_n_360, ZN => vga_com_texture_module_n_408);
  vga_com_texture_module_g16826 : AN4D0BWP7T port map(A1 => vga_com_texture_module_n_690, A2 => vga_com_texture_module_n_689, A3 => vga_com_texture_module_n_688, A4 => vga_com_texture_module_n_334, Z => vga_com_texture_module_n_407);
  vga_com_texture_module_g16827 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_361, A2 => vga_com_texture_module_n_355, B => vga_com_texture_module_n_350, ZN => vga_com_texture_module_n_406);
  vga_com_texture_module_g16828 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_frame_count(3), A2 => vga_com_texture_module_frame_count(0), B => vga_com_texture_module_n_683, ZN => vga_com_texture_module_n_405);
  vga_com_texture_module_g16829 : IOA21D1BWP7T port map(A1 => vga_com_texture_module_n_693, A2 => vga_com_texture_module_n_338, B => vga_com_texture_module_n_276, ZN => vga_com_texture_module_n_404);
  vga_com_texture_module_g16830 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_330, A2 => vga_com_texture_module_n_331, B => vga_com_texture_module_n_391, ZN => vga_com_texture_module_n_403);
  vga_com_texture_module_g16831 : IND3D0BWP7T port map(A1 => vga_com_texture_module_n_273, B1 => vga_com_texture_module_frame_count(0), B2 => vga_com_texture_module_n_366, ZN => vga_com_texture_module_n_402);
  vga_com_texture_module_g16832 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_269, A2 => vga_com_texture_module_n_364, A3 => vga_com_texture_module_n_313, ZN => vga_com_texture_module_n_416);
  vga_com_texture_module_g16833 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_283, A2 => vga_com_texture_module_n_356, A3 => vga_com_texture_module_n_350, ZN => vga_com_texture_module_n_415);
  vga_com_texture_module_g16834 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_365, A2 => vga_com_texture_module_n_356, A3 => vga_com_texture_module_n_265, ZN => vga_com_texture_module_n_413);
  vga_com_texture_module_g16835 : CKND1BWP7T port map(I => vga_com_texture_module_n_392, ZN => vga_com_texture_module_n_391);
  vga_com_texture_module_g16836 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_332, B1 => vga_com_texture_module_n_356, ZN => vga_com_texture_module_n_388);
  vga_com_texture_module_g16837 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_361, A2 => vga_com_texture_module_n_350, ZN => vga_com_texture_module_n_401);
  vga_com_texture_module_g16838 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_367, A2 => vga_com_texture_module_n_331, ZN => vga_com_texture_module_n_400);
  vga_com_texture_module_g16839 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_364, B1 => vga_com_texture_module_n_363, ZN => vga_com_texture_module_n_399);
  vga_com_texture_module_g16840 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_364, A2 => vga_com_texture_module_n_359, Z => vga_com_texture_module_n_398);
  vga_com_texture_module_g16841 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_362, B1 => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_681);
  vga_com_texture_module_g16842 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_365, A2 => vga_com_texture_module_xposition(0), Z => vga_com_texture_module_n_397);
  vga_com_texture_module_g16843 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_283, A2 => vga_com_texture_module_n_361, ZN => vga_com_texture_module_n_396);
  vga_com_texture_module_g16844 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_347, A2 => vga_com_texture_module_n_331, ZN => vga_com_texture_module_n_395);
  vga_com_texture_module_g16845 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_348, B1 => vga_com_texture_module_n_359, ZN => vga_com_texture_module_n_394);
  vga_com_texture_module_g16846 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_348, A2 => vga_com_texture_module_n_363, Z => vga_com_texture_module_n_393);
  vga_com_texture_module_g16847 : ND2D0BWP7T port map(A1 => vga_com_texture_module_n_353, A2 => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_683);
  vga_com_texture_module_g16848 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_302, A2 => vga_com_texture_module_n_349, ZN => vga_com_texture_module_n_392);
  vga_com_texture_module_g16849 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_348, A2 => vga_com_texture_module_n_314, ZN => vga_com_texture_module_n_390);
  vga_com_texture_module_g16850 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_268, A2 => vga_com_texture_module_n_345, ZN => vga_com_texture_module_n_389);
  vga_com_texture_module_g16851 : INVD1BWP7T port map(I => vga_com_texture_module_n_381, ZN => vga_com_texture_module_n_382);
  vga_com_texture_module_g16852 : INVD1BWP7T port map(I => vga_com_texture_module_n_380, ZN => vga_com_texture_module_n_379);
  vga_com_texture_module_g16853 : INVD1BWP7T port map(I => vga_com_texture_module_n_378, ZN => vga_com_texture_module_n_377);
  vga_com_texture_module_g16854 : INVD0BWP7T port map(I => vga_com_texture_module_n_376, ZN => vga_com_texture_module_n_375);
  vga_com_texture_module_g16855 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_278, A2 => vga_com_texture_module_frame_count(2), B => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_374);
  vga_com_texture_module_g16856 : OA21D0BWP7T port map(A1 => vga_com_texture_module_n_305, A2 => vga_com_texture_module_n_264, B => vga_com_texture_module_n_362, Z => vga_com_texture_module_n_373);
  vga_com_texture_module_g16857 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_682, A2 => vga_com_texture_module_n_272, A3 => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_372);
  vga_com_texture_module_g16858 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_272, A2 => vga_com_texture_module_frame_count(0), B1 => vga_com_texture_module_n_278, B2 => vga_com_texture_module_frame_count(2), ZN => vga_com_texture_module_n_371);
  vga_com_texture_module_g16859 : CKMUX2D1BWP7T port map(I0 => vga_com_bg_select(2), I1 => vga_com_texture_module_n_327, S => level_abs(0), Z => vga_com_bg_select(0));
  vga_com_texture_module_g16860 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_347, A2 => vga_com_texture_module_n_343, ZN => vga_com_texture_module_n_387);
  vga_com_texture_module_g16861 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_356, A2 => vga_com_texture_module_n_330, Z => vga_com_texture_module_n_386);
  vga_com_texture_module_g16862 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_359, A2 => vga_com_texture_module_n_330, Z => vga_com_texture_module_n_385);
  vga_com_texture_module_g16863 : AN3D1BWP7T port map(A1 => vga_com_texture_module_n_330, A2 => vga_com_texture_module_n_329, A3 => vga_com_texture_module_n_314, Z => vga_com_texture_module_n_384);
  vga_com_texture_module_g16864 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_330, A2 => vga_com_texture_module_n_329, A3 => vga_com_texture_module_n_304, ZN => vga_com_texture_module_n_383);
  vga_com_texture_module_g16865 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_274, A2 => vga_com_texture_module_n_673, B => vga_com_texture_module_n_293, ZN => vga_com_texture_module_n_370);
  vga_com_texture_module_g16866 : OA21D0BWP7T port map(A1 => vga_com_texture_module_n_669, A2 => vga_com_texture_module_n_336, B => vga_com_texture_module_n_672, Z => vga_com_texture_module_n_369);
  vga_com_texture_module_g16867 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_268, A2 => vga_com_texture_module_n_324, A3 => vga_com_texture_module_n_328, ZN => vga_com_texture_module_n_381);
  vga_com_texture_module_g16868 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_268, A2 => vga_com_texture_module_n_333, A3 => vga_com_texture_module_n_256, ZN => vga_com_texture_module_n_380);
  vga_com_texture_module_g16869 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_300, A2 => vga_com_texture_module_n_288, B1 => vga_com_texture_module_n_300, B2 => vga_com_texture_module_n_288, ZN => vga_com_texture_module_n_378);
  vga_com_texture_module_g16870 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_301, A2 => vga_com_texture_module_n_274, B1 => vga_com_texture_module_n_301, B2 => vga_com_texture_module_n_274, ZN => vga_com_texture_module_n_376);
  vga_com_texture_module_g16871 : INVD1BWP7T port map(I => vga_com_texture_module_n_358, ZN => vga_com_texture_module_n_357);
  vga_com_texture_module_g16872 : INVD1BWP7T port map(I => vga_com_texture_module_n_356, ZN => vga_com_texture_module_n_355);
  vga_com_texture_module_g16873 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_679, A2 => vga_com_texture_module_n_319, ZN => vga_com_texture_module_n_354);
  vga_com_texture_module_g16874 : NR2D0BWP7T port map(A1 => vga_com_texture_module_n_278, A2 => vga_com_texture_module_frame_count(2), ZN => vga_com_texture_module_n_353);
  vga_com_texture_module_g16875 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_320, B1 => vga_com_texture_module_n_693, ZN => vga_com_texture_module_n_368);
  vga_com_texture_module_g16876 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_322, A2 => vga_com_texture_module_yposition(1), ZN => vga_com_texture_module_n_367);
  vga_com_texture_module_g16877 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_272, B1 => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_366);
  vga_com_texture_module_g16878 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_319, B1 => vga_com_texture_module_n_679, ZN => vga_com_texture_module_n_365);
  vga_com_texture_module_g16879 : CKND2D1BWP7T port map(A1 => vga_com_texture_module_n_324, A2 => vga_com_texture_module_n_329, ZN => vga_com_texture_module_n_364);
  vga_com_texture_module_g16880 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_314, A2 => vga_com_texture_module_yposition(0), ZN => vga_com_texture_module_n_363);
  vga_com_texture_module_g16881 : IND2D0BWP7T port map(A1 => vga_com_texture_module_frame_count(0), B1 => vga_com_texture_module_n_272, ZN => vga_com_texture_module_n_362);
  vga_com_texture_module_g16882 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_335, A2 => vga_com_texture_module_xposition(0), ZN => vga_com_texture_module_n_361);
  vga_com_texture_module_g16883 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_323, A2 => vga_com_texture_module_yposition(0), Z => vga_com_texture_module_n_360);
  vga_com_texture_module_g16884 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_313, A2 => vga_com_texture_module_yposition(0), ZN => vga_com_texture_module_n_359);
  vga_com_texture_module_g16885 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_332, A2 => vga_com_texture_module_yposition(0), ZN => vga_com_texture_module_n_358);
  vga_com_texture_module_g16886 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_323, B1 => vga_com_texture_module_yposition(0), ZN => vga_com_texture_module_n_356);
  vga_com_texture_module_g16887 : INVD0BWP7T port map(I => vga_com_texture_module_n_345, ZN => vga_com_texture_module_n_344);
  vga_com_texture_module_g16888 : INVD1BWP7T port map(I => vga_com_texture_module_n_343, ZN => vga_com_texture_module_n_342);
  vga_com_texture_module_g16889 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_285, A2 => vga_com_texture_module_n_263, B1 => vga_com_texture_module_n_305, B2 => vga_com_texture_module_frame_count(2), ZN => vga_com_texture_module_n_341);
  vga_com_texture_module_g16890 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_291, A2 => vga_com_texture_module_n_286, B => vga_com_texture_module_n_318, ZN => vga_com_texture_module_n_340);
  vga_com_texture_module_g16891 : OAI221D0BWP7T port map(A1 => vga_com_texture_module_n_264, A2 => vga_com_texture_module_frame_count(1), B1 => vga_com_texture_module_n_260, B2 => vga_com_texture_module_frame_count(2), C => vga_com_texture_module_frame_count(0), ZN => vga_com_texture_module_n_339);
  vga_com_texture_module_g16892 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_277, A2 => vga_com_texture_module_n_306, B => vga_com_texture_module_n_320, ZN => vga_com_texture_module_n_338);
  vga_com_texture_module_g16893 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_277, A2 => vga_com_texture_module_n_308, B => vga_com_texture_module_n_320, ZN => vga_com_texture_module_n_337);
  vga_com_texture_module_g16894 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_299, A2 => vga_com_texture_module_n_290, B => vga_com_texture_module_n_303, ZN => vga_com_texture_module_n_352);
  vga_com_texture_module_g16895 : AOI32D1BWP7T port map(A1 => vga_com_texture_module_n_270, A2 => vga_com_texture_module_n_279, A3 => vga_com_texture_module_xposition(3), B1 => vga_com_texture_module_n_271, B2 => vga_com_texture_module_n_298, ZN => vga_com_texture_module_n_351);
  vga_com_texture_module_g16896 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_298, A2 => vga_com_texture_module_n_265, A3 => vga_com_texture_module_xposition(1), ZN => vga_com_texture_module_n_350);
  vga_com_texture_module_g16897 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_296, A2 => vga_com_texture_module_n_265, A3 => vga_com_texture_module_n_256, ZN => vga_com_texture_module_n_349);
  vga_com_texture_module_g16898 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_269, A2 => vga_com_texture_module_n_309, A3 => vga_com_texture_module_n_270, ZN => vga_com_texture_module_n_348);
  vga_com_texture_module_g16899 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_302, A2 => vga_com_texture_module_n_316, ZN => vga_com_texture_module_n_347);
  vga_com_texture_module_g16900 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_304, B1 => vga_com_texture_module_yposition(1), B2 => vga_com_texture_module_n_21, ZN => vga_com_texture_module_n_346);
  vga_com_texture_module_g16901 : AOI31D0BWP7T port map(A1 => vga_com_texture_module_n_271, A2 => vga_com_texture_module_xposition(2), A3 => vga_com_texture_module_xposition(3), B => vga_com_texture_module_xposition(4), ZN => vga_com_texture_module_n_345);
  vga_com_texture_module_g16902 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_28, A2 => vga_com_texture_module_n_316, ZN => vga_com_texture_module_n_343);
  vga_com_texture_module_g16903 : INVD1BWP7T port map(I => vga_com_texture_module_n_288, ZN => vga_com_texture_module_n_336);
  vga_com_texture_module_g16904 : INVD0BWP7T port map(I => vga_com_texture_module_n_293, ZN => vga_com_texture_module_n_674);
  vga_com_texture_module_g16905 : INVD1BWP7T port map(I => vga_com_texture_module_n_328, ZN => vga_com_texture_module_n_329);
  vga_com_texture_module_g16906 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_297, A2 => level_abs(1), ZN => vga_com_texture_module_n_327);
  vga_com_texture_module_g16907 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_308, B1 => vga_com_texture_module_n_691, ZN => vga_com_texture_module_n_326);
  vga_com_texture_module_g16908 : IND2D1BWP7T port map(A1 => level_abs(0), B1 => vga_com_texture_module_n_297, ZN => vga_com_bg_select(1));
  vga_com_texture_module_g16909 : IND2D1BWP7T port map(A1 => level_abs(1), B1 => vga_com_texture_module_n_297, ZN => vga_com_bg_select(2));
  vga_com_texture_module_g16910 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_298, A2 => vga_com_texture_module_n_256, Z => vga_com_texture_module_n_335);
  vga_com_texture_module_g16911 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_687, B1 => vga_com_texture_module_n_306, ZN => vga_com_texture_module_n_334);
  vga_com_texture_module_g16912 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_309, A2 => vga_com_texture_module_n_265, ZN => vga_com_texture_module_n_333);
  vga_com_texture_module_g16913 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_304, A2 => vga_com_texture_module_yposition(1), ZN => vga_com_texture_module_n_332);
  vga_com_texture_module_g16914 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_299, A2 => vga_com_texture_module_n_286, ZN => vga_com_texture_module_n_331);
  vga_com_texture_module_g16915 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_307, A2 => vga_com_texture_module_n_21, Z => vga_com_texture_module_n_330);
  vga_com_texture_module_g16916 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_307, A2 => FE_PHN253_vga_com_texture_module_yposition_0, ZN => vga_com_texture_module_n_328);
  vga_com_texture_module_g16917 : INVD0BWP7T port map(I => vga_com_texture_module_n_322, ZN => vga_com_texture_module_n_321);
  vga_com_texture_module_g16918 : INVD0BWP7T port map(I => vga_com_texture_module_n_317, ZN => vga_com_texture_module_n_318);
  vga_com_texture_module_g16919 : INVD0BWP7T port map(I => vga_com_texture_module_n_316, ZN => vga_com_texture_module_n_315);
  vga_com_texture_module_g16920 : INVD1BWP7T port map(I => vga_com_texture_module_n_314, ZN => vga_com_texture_module_n_313);
  vga_com_texture_module_g16921 : AO31D1BWP7T port map(A1 => vga_com_texture_module_n_280, A2 => vga_com_vcount(5), A3 => FE_PHN239_vga_com_vcount_8, B => FE_PHN241_vga_com_vcount_9, Z => vga_done);
  vga_com_texture_module_g16922 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_285, A2 => vga_com_texture_module_frame_count(2), B => vga_com_texture_module_n_305, ZN => vga_com_texture_module_n_312);
  vga_com_texture_module_g16923 : IAO21D0BWP7T port map(A1 => vga_com_texture_module_n_285, A2 => vga_com_texture_module_n_264, B => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_311);
  vga_com_texture_module_g16924 : INR2D0BWP7T port map(A1 => vga_com_texture_module_n_305, B1 => vga_com_texture_module_n_273, ZN => vga_com_texture_module_n_325);
  vga_com_texture_module_g16925 : AN3D1BWP7T port map(A1 => vga_com_texture_module_n_271, A2 => vga_com_texture_module_n_279, A3 => vga_com_texture_module_xposition(3), Z => vga_com_texture_module_n_324);
  vga_com_texture_module_g16926 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_290, A2 => vga_com_texture_module_n_25, A3 => vga_com_texture_module_yposition(1), ZN => vga_com_texture_module_n_323);
  vga_com_texture_module_g16927 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_304, A2 => vga_com_texture_module_n_21, ZN => vga_com_texture_module_n_322);
  vga_com_texture_module_g16928 : OAI31D0BWP7T port map(A1 => vga_com_texture_module_n_688, A2 => vga_com_texture_module_n_689, A3 => vga_com_texture_module_n_690, B => vga_com_texture_module_n_691, ZN => vga_com_texture_module_n_320);
  vga_com_texture_module_g16929 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_296, A2 => vga_com_texture_module_xposition(1), ZN => vga_com_texture_module_n_319);
  vga_com_texture_module_g16930 : IND2D1BWP7T port map(A1 => vga_com_texture_module_yposition(4), B1 => vga_com_texture_module_n_299, ZN => vga_com_texture_module_n_317);
  vga_com_texture_module_g16931 : CKND2D1BWP7T port map(A1 => vga_com_texture_module_n_310, A2 => vga_com_texture_module_n_271, ZN => vga_com_texture_module_n_316);
  vga_com_texture_module_g16932 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_286, A2 => vga_com_texture_module_n_25, A3 => vga_com_texture_module_yposition(1), ZN => vga_com_texture_module_n_314);
  vga_com_texture_module_g16933 : INVD0BWP7T port map(I => vga_com_texture_module_n_304, ZN => vga_com_texture_module_n_303);
  vga_com_texture_module_g16934 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_281, B1 => vga_com_texture_module_xposition(4), ZN => vga_com_texture_module_n_310);
  vga_com_texture_module_g16935 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_281, A2 => vga_com_texture_module_xposition(4), ZN => vga_com_texture_module_n_309);
  vga_com_texture_module_g16936 : INR2XD0BWP7T port map(A1 => vga_com_texture_module_n_292, B1 => vga_com_texture_module_n_686, ZN => vga_com_texture_module_n_308);
  vga_com_texture_module_g16937 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_712, B1 => vga_com_texture_module_frame_count(2), ZN => vga_com_texture_module_n_676);
  vga_com_texture_module_g16938 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_291, B1 => vga_com_texture_module_n_290, ZN => vga_com_texture_module_n_307);
  vga_com_texture_module_g16939 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_292, B1 => vga_com_texture_module_n_686, ZN => vga_com_texture_module_n_306);
  vga_com_texture_module_g16940 : ND2D0BWP7T port map(A1 => vga_com_texture_module_n_712, A2 => vga_com_texture_module_n_263, ZN => vga_com_texture_module_n_305);
  vga_com_texture_module_g16941 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_286, A2 => vga_com_texture_module_yposition(3), ZN => vga_com_texture_module_n_304);
  vga_com_texture_module_g16942 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_678, A2 => vga_com_texture_module_n_289, ZN => vga_com_texture_module_n_302);
  vga_com_texture_module_g16943 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_yposition(1), A2 => yplayer(1), B1 => vga_com_texture_module_yposition(1), B2 => yplayer(1), ZN => vga_com_texture_module_n_301);
  vga_com_texture_module_g16944 : MAOI22D0BWP7T port map(A1 => xplayer(1), A2 => vga_com_texture_module_xposition(1), B1 => xplayer(1), B2 => vga_com_texture_module_xposition(1), ZN => vga_com_texture_module_n_300);
  vga_com_texture_module_g16945 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_260, A2 => vga_com_texture_module_frame_count(0), B => vga_com_texture_module_n_278, ZN => vga_com_texture_module_n_682);
  vga_com_texture_module_g16946 : NR3D0BWP7T port map(A1 => vga_com_texture_module_yposition(0), A2 => vga_com_texture_module_n_25, A3 => vga_com_texture_module_yposition(1), ZN => vga_com_texture_module_n_299);
  vga_com_texture_module_g16947 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_257, A2 => vga_com_texture_module_xposition(2), A3 => vga_com_texture_module_xposition(4), ZN => vga_com_texture_module_n_298);
  vga_com_texture_module_g16948 : NR3D0BWP7T port map(A1 => level_abs(2), A2 => level_abs(4), A3 => level_abs(3), ZN => vga_com_texture_module_n_297);
  vga_com_texture_module_g16949 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_279, B1 => vga_com_texture_module_xposition(3), ZN => vga_com_texture_module_n_296);
  vga_com_texture_module_g16950 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_xposition(0), A2 => xplayer(0), B1 => xplayer(0), B2 => vga_com_texture_module_xposition(0), ZN => vga_com_texture_module_n_295);
  vga_com_texture_module_g16951 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_yposition(0), A2 => yplayer(0), B1 => yplayer(0), B2 => vga_com_texture_module_yposition(0), ZN => vga_com_texture_module_n_294);
  vga_com_texture_module_g16952 : INVD0BWP7T port map(I => vga_com_texture_module_n_679, ZN => vga_com_texture_module_n_28);
  vga_com_texture_module_g16953 : INVD1BWP7T port map(I => vga_com_texture_module_n_283, ZN => vga_com_texture_module_n_678);
  vga_com_texture_module_g16954 : ND2D1BWP7T port map(A1 => xplayer(3), A2 => vga_com_texture_module_n_257, ZN => vga_com_texture_module_n_282);
  vga_com_texture_module_g16955 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_266, A2 => yplayer(1), ZN => vga_com_texture_module_n_673);
  vga_com_texture_module_g16956 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_266, A2 => yplayer(1), ZN => vga_com_texture_module_n_293);
  vga_com_texture_module_g16957 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_684, A2 => vga_com_texture_module_n_685, ZN => vga_com_texture_module_n_292);
  vga_com_texture_module_g16958 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_266, A2 => vga_com_texture_module_n_25, ZN => vga_com_texture_module_n_291);
  vga_com_texture_module_g16959 : INR2D1BWP7T port map(A1 => xplayer(1), B1 => vga_com_texture_module_xposition(1), ZN => vga_com_texture_module_n_669);
  vga_com_texture_module_g16960 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_7, A2 => vga_com_texture_module_yposition(4), ZN => vga_com_texture_module_n_290);
  vga_com_texture_module_g16961 : NR2D1BWP7T port map(A1 => game_state(0), A2 => game_state(1), ZN => vga_com_texture_module_n_289);
  vga_com_texture_module_g16962 : CKND2D1BWP7T port map(A1 => vga_com_texture_module_n_265, A2 => xplayer(0), ZN => vga_com_texture_module_n_288);
  vga_com_texture_module_g16963 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_697, A2 => vga_com_texture_module_n_696, ZN => vga_com_texture_module_n_287);
  vga_com_texture_module_g16964 : NR2D1BWP7T port map(A1 => vga_com_texture_module_yposition(2), A2 => vga_com_texture_module_yposition(4), ZN => vga_com_texture_module_n_286);
  vga_com_texture_module_g16965 : NR2D0BWP7T port map(A1 => vga_com_texture_module_frame_count(0), A2 => vga_com_texture_module_frame_count(1), ZN => vga_com_texture_module_n_285);
  vga_com_texture_module_g16966 : INR2D1BWP7T port map(A1 => game_state(1), B1 => game_state(0), ZN => vga_com_texture_module_n_679);
  vga_com_texture_module_g16967 : ND2D1BWP7T port map(A1 => game_state(0), A2 => game_state(1), ZN => vga_com_texture_module_n_283);
  vga_com_texture_module_g16968 : CKND1BWP7T port map(I => vga_com_texture_module_n_667, ZN => vga_com_texture_module_n_280);
  vga_com_texture_module_g16969 : INVD1BWP7T port map(I => vga_com_texture_module_n_276, ZN => vga_com_texture_module_n_275);
  vga_com_texture_module_g16970 : INVD1BWP7T port map(I => vga_com_texture_module_n_271, ZN => vga_com_texture_module_n_270);
  vga_com_texture_module_g16971 : INVD1BWP7T port map(I => vga_com_texture_module_n_269, ZN => vga_com_texture_module_n_268);
  vga_com_texture_module_g16972 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_257, A2 => xplayer(3), ZN => vga_com_texture_module_n_267);
  vga_com_texture_module_g16973 : NR2D0BWP7T port map(A1 => vga_com_texture_module_xposition(2), A2 => vga_com_texture_module_xposition(3), ZN => vga_com_texture_module_n_281);
  vga_com_texture_module_g16974 : IND2D1BWP7T port map(A1 => xplayer(1), B1 => vga_com_texture_module_xposition(1), ZN => vga_com_texture_module_n_672);
  vga_com_texture_module_g16975 : ND2D1BWP7T port map(A1 => vga_com_vcount(6), A2 => FE_PHN238_vga_com_vcount_7, ZN => vga_com_texture_module_n_667);
  vga_com_texture_module_g16976 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_259, A2 => vga_com_texture_module_xposition(4), ZN => vga_com_texture_module_n_279);
  vga_com_texture_module_g16977 : ND2D0BWP7T port map(A1 => vga_com_texture_module_n_260, A2 => vga_com_texture_module_frame_count(0), ZN => vga_com_texture_module_n_278);
  vga_com_texture_module_g16978 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_691, A2 => vga_com_texture_module_n_687, ZN => vga_com_texture_module_n_277);
  vga_com_texture_module_g16979 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_693, A2 => vga_com_texture_module_n_692, ZN => vga_com_texture_module_n_276);
  vga_com_texture_module_g16980 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_21, A2 => yplayer(0), ZN => vga_com_texture_module_n_274);
  vga_com_texture_module_g16981 : NR2D0BWP7T port map(A1 => vga_com_texture_module_frame_count(2), A2 => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_273);
  vga_com_texture_module_g16982 : ND2D0BWP7T port map(A1 => vga_com_texture_module_frame_count(0), A2 => vga_com_texture_module_frame_count(1), ZN => vga_com_texture_module_n_712);
  vga_com_texture_module_g16983 : NR2D0BWP7T port map(A1 => vga_com_texture_module_frame_count(2), A2 => vga_com_texture_module_frame_count(1), ZN => vga_com_texture_module_n_272);
  vga_com_texture_module_g16984 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_265, A2 => vga_com_texture_module_n_256, ZN => vga_com_texture_module_n_271);
  vga_com_texture_module_g16985 : IND2D1BWP7T port map(A1 => game_state(1), B1 => game_state(0), ZN => vga_com_texture_module_n_269);
  vga_com_texture_module_g16990 : INVD0BWP7T port map(I => vga_com_texture_module_n_693, ZN => vga_com_texture_module_n_262);
  vga_com_texture_module_column_reg_0 : DFQD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_188, Q => vga_com_column(0));
  vga_com_texture_module_frame_count_reg_0 : DFCNQD1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_com_texture_module_timer1(4), D => vga_com_texture_module_n_71, Q => vga_com_texture_module_frame_count(0));
  vga_com_texture_module_hcount_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN352_vga_com_texture_module_n_52, CP => CTS_23, D => vga_com_texture_module_n_139, Q => vga_com_hcount(1));
  vga_com_texture_module_hcount_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN203_vga_com_texture_module_n_79, CP => CTS_23, D => vga_com_texture_module_n_139, Q => vga_com_hcount(2));
  vga_com_texture_module_hcount_reg_3 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_105, CP => CTS_23, D => vga_com_texture_module_n_139, Q => vga_com_hcount(3));
  vga_com_texture_module_hcount_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN216_vga_com_texture_module_n_115, CP => CTS_23, D => vga_com_texture_module_n_139, Q => vga_com_hcount(4));
  vga_com_texture_module_hcount_reg_7 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_139, CP => CTS_23, D => vga_com_texture_module_n_217, Q => vga_com_hcount(7));
  vga_com_texture_module_hcount_reg_9 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_139, CP => CTS_23, D => vga_com_texture_module_n_245, Q => vga_com_hcount(9));
  vga_com_texture_module_hvis_reg_3 : DFXQD1BWP7T port map(CP => CTS_23, DA => FE_PHN362_vga_com_texture_module_n_176, DB => vga_com_texture_module_n_165, Q => vga_com_texture_module_hvis(3), SA => FE_PHN370_vga_com_texture_module_hvis_3);
  vga_com_texture_module_hvis_reg_6 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN353_vga_com_texture_module_n_174, Q => vga_com_texture_module_hvis(6));
  vga_com_texture_module_row_reg_0 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_151, CP => CTS_23, D => vga_com_texture_module_n_154, Q => vga_com_row(0));
  vga_com_texture_module_row_reg_1 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_191, CP => CTS_23, D => vga_com_texture_module_n_154, Q => vga_com_row(1));
  vga_com_texture_module_row_reg_2 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_154, CP => CTS_23, D => vga_com_texture_module_n_228, Q => vga_com_row(2));
  vga_com_texture_module_timer1_reg_1 : EDFCND1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_done, D => vga_com_texture_module_timer1(1), E => vga_com_texture_module_timer1(0), Q => UNCONNECTED, QN => vga_com_texture_module_timer1(1));
  vga_com_texture_module_timer1_reg_2 : DFCNQD1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_done, D => vga_com_texture_module_n_82, Q => vga_com_texture_module_timer1(2));
  vga_com_texture_module_timer1_reg_3 : DFCNQD1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_done, D => vga_com_texture_module_n_103, Q => vga_com_texture_module_timer1(3));
  vga_com_texture_module_timer1_reg_5 : DFCNQD1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_done, D => vga_com_texture_module_n_138, Q => vga_com_timer1(5));
  vga_com_texture_module_vcount_reg_1 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN311_vga_com_texture_module_n_201, Q => vga_com_vcount(1));
  vga_com_texture_module_vcount_reg_2 : DFXQD1BWP7T port map(CP => CTS_23, DA => vga_com_texture_module_n_210, DB => FE_PHN408_vga_com_texture_module_n_193, Q => FE_PHN401_vga_com_vcount_2, SA => FE_PHN231_vga_com_vcount_2);
  vga_com_texture_module_vcount_reg_3 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN312_vga_com_texture_module_n_242, Q => vga_com_vcount(3));
  vga_com_texture_module_vcount_reg_4 : DFQD0BWP7T port map(CP => CTS_23, D => FE_PHN344_vga_com_texture_module_n_240, Q => vga_com_vcount(4));
  vga_com_texture_module_vvis_reg_1 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN358_vga_com_texture_module_n_238, Q => vga_com_texture_module_vvis(1));
  vga_com_texture_module_vvis_reg_3 : DFQD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_248, Q => vga_com_texture_module_vvis(3));
  vga_com_texture_module_vvis_reg_5 : DFQD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_253, Q => vga_com_texture_module_vvis(5));
  vga_com_texture_module_vvis_reg_6 : DFQD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_241, Q => vga_com_texture_module_vvis(6));
  vga_com_texture_module_xposition_reg_4 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_136, CP => CTS_23, D => FE_PHN354_vga_com_texture_module_n_239, Q => FE_PHN254_vga_com_texture_module_xposition_4);
  vga_com_texture_module_yposition_reg_4 : DFKCNQD1BWP7T port map(CN => vga_com_texture_module_n_146, CP => CTS_23, D => vga_com_texture_module_n_254, Q => vga_com_texture_module_yposition(4));
  vga_com_texture_module_g11162 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_250, A2 => vga_com_texture_module_yposition(4), B1 => vga_com_texture_module_n_250, B2 => vga_com_texture_module_yposition(4), ZN => FE_PHN342_vga_com_texture_module_n_254);
  vga_com_texture_module_g11171 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_246, A2 => vga_com_texture_module_n_199, ZN => FE_PHN327_vga_com_texture_module_n_253);
  vga_com_texture_module_g11172 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_225, A2 => vga_com_texture_module_yposition(3), B1 => vga_com_texture_module_n_225, B2 => vga_com_texture_module_yposition(3), ZN => FE_PHN404_vga_com_texture_module_n_252);
  vga_com_texture_module_g11173 : AO22D0BWP7T port map(A1 => vga_com_texture_module_n_243, A2 => FE_PHN241_vga_com_vcount_9, B1 => FE_PHN239_vga_com_vcount_8, B2 => vga_com_texture_module_n_219, Z => vga_com_texture_module_n_251);
  vga_com_texture_module_g11177 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_225, B1 => vga_com_texture_module_yposition(3), ZN => vga_com_texture_module_n_250);
  vga_com_texture_module_g11183 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_234, A2 => vga_com_texture_module_n_194, A3 => vga_com_texture_module_n_152, ZN => vga_com_texture_module_n_249);
  vga_com_texture_module_g11184 : OAI211D1BWP7T port map(A1 => vga_com_texture_module_vvis(3), A2 => vga_com_texture_module_n_205, B => vga_com_texture_module_n_236, C => vga_com_texture_module_n_152, ZN => FE_PHN318_vga_com_texture_module_n_248);
  vga_com_texture_module_g11185 : OAI221D0BWP7T port map(A1 => vga_com_texture_module_n_227, A2 => vga_com_texture_module_n_9, B1 => vga_com_texture_module_vvis(4), B2 => vga_com_texture_module_n_215, C => vga_com_texture_module_n_152, ZN => vga_com_texture_module_n_247);
  vga_com_texture_module_g11186 : AOI222D0BWP7T port map(A1 => vga_com_texture_module_n_230, A2 => vga_com_texture_module_vvis(5), B1 => vga_com_texture_module_n_214, B2 => vga_com_texture_module_vvis(4), C1 => vga_com_texture_module_n_153, C2 => yplayer(0), ZN => vga_com_texture_module_n_246);
  vga_com_texture_module_g11187 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_220, A2 => vga_com_hcount(8), B => FE_PHN235_vga_com_hcount_9, Z => vga_com_texture_module_n_245);
  vga_com_texture_module_g11188 : AO32D1BWP7T port map(A1 => vga_com_texture_module_n_192, A2 => vga_com_texture_module_n_10, A3 => vga_com_vcount(6), B1 => vga_com_texture_module_n_233, B2 => FE_PHN238_vga_com_vcount_7, Z => vga_com_texture_module_n_244);
  vga_com_texture_module_g11193 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_178, A2 => vga_com_texture_module_n_4, B => vga_com_texture_module_n_235, Z => vga_com_texture_module_n_243);
  vga_com_texture_module_g11194 : IOA21D1BWP7T port map(A1 => vga_com_texture_module_n_221, A2 => vga_com_vcount(3), B => vga_com_texture_module_n_224, ZN => vga_com_texture_module_n_242);
  vga_com_texture_module_g11195 : OAI221D0BWP7T port map(A1 => vga_com_texture_module_n_203, A2 => FE_PHN101_vga_com_texture_module_vvis_6, B1 => vga_com_texture_module_n_50, B2 => vga_com_texture_module_n_152, C => vga_com_texture_module_n_237, ZN => vga_com_texture_module_n_241);
  vga_com_texture_module_g11196 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_212, A2 => vga_com_vcount(4), B1 => vga_com_texture_module_n_222, B2 => vga_com_vcount(4), ZN => vga_com_texture_module_n_240);
  vga_com_texture_module_g11197 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_195, A2 => vga_com_texture_module_xposition(4), B1 => vga_com_texture_module_n_195, B2 => vga_com_texture_module_xposition(4), ZN => vga_com_texture_module_n_239);
  vga_com_texture_module_g11198 : OAI211D1BWP7T port map(A1 => vga_com_texture_module_n_54, A2 => vga_com_texture_module_n_180, B => vga_com_texture_module_n_207, C => vga_com_texture_module_n_152, ZN => vga_com_texture_module_n_238);
  vga_com_texture_module_g11199 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_208, A2 => vga_com_texture_module_n_136, B => FE_PHN101_vga_com_texture_module_vvis_6, ZN => vga_com_texture_module_n_237);
  vga_com_texture_module_g11200 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_218, A2 => vga_com_texture_module_n_200, B => vga_com_texture_module_vvis(3), ZN => vga_com_texture_module_n_236);
  vga_com_texture_module_g11205 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_218, A2 => vga_com_texture_module_vvis(2), B1 => vga_com_texture_module_n_180, B2 => vga_com_texture_module_n_81, ZN => vga_com_texture_module_n_234);
  vga_com_texture_module_g11206 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_178, A2 => vga_com_texture_module_n_2, B => vga_com_texture_module_n_226, Z => vga_com_texture_module_n_233);
  vga_com_texture_module_g11207 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_220, A2 => vga_com_texture_module_n_1, B1 => vga_com_texture_module_n_220, B2 => vga_com_texture_module_n_1, ZN => FE_PHN343_vga_com_texture_module_n_232);
  vga_com_texture_module_g11208 : OAI32D1BWP7T port map(A1 => vga_com_vcount(5), A2 => vga_com_texture_module_n_85, A3 => vga_com_texture_module_n_177, B1 => FE_PHN217_vga_com_texture_module_n_6, B2 => vga_com_texture_module_n_211, ZN => vga_com_texture_module_n_231);
  vga_com_texture_module_g11209 : OAI221D0BWP7T port map(A1 => vga_com_texture_module_n_180, A2 => vga_com_texture_module_vvis(4), B1 => vga_com_texture_module_n_9, B2 => vga_com_texture_module_n_182, C => vga_com_texture_module_n_227, ZN => vga_com_texture_module_n_230);
  vga_com_texture_module_g11210 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_183, A2 => vga_com_texture_module_yposition(2), B1 => vga_com_texture_module_n_183, B2 => vga_com_texture_module_yposition(2), ZN => vga_com_texture_module_n_229);
  vga_com_texture_module_g11211 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_184, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_texture_module_n_184, B2 => FE_OFN4_vga_com_row_2, ZN => vga_com_texture_module_n_228);
  vga_com_texture_module_g11212 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_178, A2 => vga_com_texture_module_n_667, B => vga_com_texture_module_n_226, Z => vga_com_texture_module_n_235);
  vga_com_texture_module_g11220 : IND3D1BWP7T port map(A1 => vga_com_vcount(3), B1 => FE_PHN231_vga_com_vcount_2, B2 => vga_com_texture_module_n_193, ZN => vga_com_texture_module_n_224);
  vga_com_texture_module_g11221 : OAI211D1BWP7T port map(A1 => xplayer(0), A2 => vga_com_texture_module_n_120, B => vga_com_texture_module_n_189, C => vga_com_texture_module_n_197, ZN => FE_PHN300_vga_com_texture_module_n_223);
  vga_com_texture_module_g11222 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_178, A2 => vga_com_texture_module_n_32, B => vga_com_texture_module_n_210, Z => vga_com_texture_module_n_222);
  vga_com_texture_module_g11223 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_177, A2 => FE_PHN231_vga_com_vcount_2, B => vga_com_texture_module_n_209, ZN => vga_com_texture_module_n_221);
  vga_com_texture_module_g11224 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_179, A2 => vga_com_texture_module_n_100, B => vga_com_texture_module_n_218, C => vga_com_texture_module_n_196, ZN => vga_com_texture_module_n_227);
  vga_com_texture_module_g11225 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_177, A2 => vga_com_vcount(5), B => vga_com_texture_module_n_211, ZN => vga_com_texture_module_n_226);
  vga_com_texture_module_g11226 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_183, B1 => vga_com_texture_module_yposition(2), ZN => vga_com_texture_module_n_225);
  vga_com_texture_module_g11227 : HA1D0BWP7T port map(A => FE_PHN161_vga_com_hcount_7, B => vga_com_texture_module_n_170, CO => vga_com_texture_module_n_220, S => vga_com_texture_module_n_217);
  vga_com_texture_module_g11228 : AO211D0BWP7T port map(A1 => vga_com_texture_module_n_168, A2 => vga_com_texture_module_hvis(2), B => vga_com_texture_module_n_155, C => vga_com_texture_module_n_149, Z => FE_PHN341_vga_com_texture_module_n_216);
  vga_com_texture_module_g11229 : IAO21D0BWP7T port map(A1 => vga_com_texture_module_n_182, A2 => vga_com_texture_module_n_78, B => vga_com_texture_module_n_198, ZN => vga_com_texture_module_n_215);
  vga_com_texture_module_g11230 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_198, B1 => vga_com_texture_module_vvis(5), ZN => vga_com_texture_module_n_214);
  vga_com_texture_module_g11231 : AO221D0BWP7T port map(A1 => vga_com_texture_module_n_167, A2 => vga_com_texture_module_n_16, B1 => vga_com_texture_module_n_136, B2 => FE_PHN391_vga_com_texture_module_vvis_0, C => vga_com_texture_module_n_153, Z => vga_com_texture_module_n_213);
  vga_com_texture_module_g11232 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_32, B1 => vga_com_texture_module_n_193, ZN => vga_com_texture_module_n_212);
  vga_com_texture_module_g11233 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_192, B1 => vga_com_texture_module_n_667, ZN => vga_com_texture_module_n_219);
  vga_com_texture_module_g11234 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_182, A2 => vga_com_texture_module_n_42, B => vga_com_texture_module_n_135, ZN => vga_com_texture_module_n_218);
  vga_com_texture_module_g11238 : INVD1BWP7T port map(I => vga_com_texture_module_n_209, ZN => vga_com_texture_module_n_210);
  vga_com_texture_module_g11239 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_182, A2 => vga_com_texture_module_n_90, B1 => vga_com_texture_module_n_180, B2 => vga_com_texture_module_n_106, ZN => vga_com_texture_module_n_208);
  vga_com_texture_module_g11240 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_181, A2 => vga_com_texture_module_n_54, B1 => vga_com_texture_module_n_136, B2 => vga_com_texture_module_vvis(1), ZN => vga_com_texture_module_n_207);
  vga_com_texture_module_g11241 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_186, A2 => FE_PHN17_vga_com_texture_module_n_20, B => vga_com_texture_module_n_175, ZN => vga_com_texture_module_n_206);
  vga_com_texture_module_g11242 : OA21D0BWP7T port map(A1 => vga_com_texture_module_n_180, A2 => vga_com_texture_module_n_94, B => vga_com_texture_module_n_194, Z => vga_com_texture_module_n_205);
  vga_com_texture_module_g11243 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_159, A2 => vga_com_texture_module_xposition(3), B1 => vga_com_texture_module_n_159, B2 => vga_com_texture_module_xposition(3), ZN => vga_com_texture_module_n_204);
  vga_com_texture_module_g11244 : OA21D0BWP7T port map(A1 => vga_com_texture_module_n_180, A2 => vga_com_texture_module_n_107, B => vga_com_texture_module_n_199, Z => vga_com_texture_module_n_203);
  vga_com_texture_module_g11245 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_158, A2 => vga_com_texture_module_n_62, B1 => vga_com_texture_module_n_185, B2 => vga_com_column(2), ZN => vga_com_texture_module_n_202);
  vga_com_texture_module_g11246 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_177, A2 => vga_com_texture_module_n_49, B1 => vga_com_texture_module_n_166, B2 => vga_com_vcount(1), ZN => vga_com_texture_module_n_201);
  vga_com_texture_module_g11247 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_180, A2 => vga_com_texture_module_n_75, B1 => vga_com_texture_module_n_182, B2 => vga_com_texture_module_n_8, ZN => vga_com_texture_module_n_200);
  vga_com_texture_module_g11248 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_178, A2 => vga_com_texture_module_n_85, B => vga_com_texture_module_n_166, ZN => vga_com_texture_module_n_211);
  vga_com_texture_module_g11249 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_178, A2 => vga_com_texture_module_n_33, B => vga_com_texture_module_n_166, ZN => vga_com_texture_module_n_209);
  vga_com_texture_module_g11250 : IOA21D1BWP7T port map(A1 => vga_com_texture_module_n_169, A2 => vga_com_texture_module_n_161, B => vga_com_texture_module_hvis(5), ZN => vga_com_texture_module_n_197);
  vga_com_texture_module_g11251 : NR2D0BWP7T port map(A1 => vga_com_texture_module_n_182, A2 => vga_com_texture_module_n_668, ZN => vga_com_texture_module_n_196);
  vga_com_texture_module_g11252 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_181, A2 => vga_com_texture_module_n_90, ZN => vga_com_texture_module_n_199);
  vga_com_texture_module_g11253 : NR2D0BWP7T port map(A1 => vga_com_texture_module_n_180, A2 => vga_com_texture_module_n_100, ZN => vga_com_texture_module_n_198);
  vga_com_texture_module_g11258 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_147, A2 => FE_OFN3_vga_com_row_1, B1 => vga_com_texture_module_n_147, B2 => FE_OFN3_vga_com_row_1, ZN => vga_com_texture_module_n_191);
  vga_com_texture_module_g11259 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_148, A2 => vga_com_texture_module_yposition(1), B1 => vga_com_texture_module_n_148, B2 => vga_com_texture_module_yposition(1), ZN => vga_com_texture_module_n_190);
  vga_com_texture_module_g11260 : AOI32D1BWP7T port map(A1 => vga_com_texture_module_n_160, A2 => vga_com_texture_module_n_22, A3 => vga_com_texture_module_hvis(4), B1 => vga_com_texture_module_n_144, B2 => vga_com_texture_module_n_89, ZN => vga_com_texture_module_n_189);
  vga_com_texture_module_g11261 : IOA21D1BWP7T port map(A1 => vga_com_texture_module_n_173, A2 => vga_com_column(0), B => vga_com_texture_module_n_172, ZN => vga_com_texture_module_n_188);
  vga_com_texture_module_g11262 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_163, A2 => vga_com_texture_module_hvis(4), B1 => vga_com_texture_module_n_169, B2 => vga_com_texture_module_n_5, ZN => FE_PHN309_vga_com_texture_module_n_187);
  vga_com_texture_module_g11263 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_159, B1 => vga_com_texture_module_xposition(3), ZN => vga_com_texture_module_n_195);
  vga_com_texture_module_g11264 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_181, A2 => vga_com_texture_module_n_42, A3 => vga_com_texture_module_n_8, ZN => vga_com_texture_module_n_194);
  vga_com_texture_module_g11265 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_177, A2 => vga_com_texture_module_n_33, ZN => vga_com_texture_module_n_193);
  vga_com_texture_module_g11266 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_177, A2 => vga_com_texture_module_n_85, A3 => FE_PHN217_vga_com_texture_module_n_6, ZN => vga_com_texture_module_n_192);
  vga_com_texture_module_g11267 : INVD0BWP7T port map(I => vga_com_texture_module_n_185, ZN => vga_com_texture_module_n_186);
  vga_com_texture_module_g11268 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_173, B1 => vga_com_texture_module_n_172, ZN => vga_com_texture_module_n_185);
  vga_com_texture_module_g11269 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_147, B1 => FE_OFN3_vga_com_row_1, ZN => vga_com_texture_module_n_184);
  vga_com_texture_module_g11270 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_148, B1 => vga_com_texture_module_yposition(1), ZN => vga_com_texture_module_n_183);
  vga_com_texture_module_g11273 : INVD0BWP7T port map(I => vga_com_texture_module_n_182, ZN => vga_com_texture_module_n_181);
  vga_com_texture_module_g11274 : INVD0BWP7T port map(I => vga_com_texture_module_n_180, ZN => vga_com_texture_module_n_179);
  vga_com_texture_module_g11275 : INVD1BWP7T port map(I => vga_com_texture_module_n_178, ZN => vga_com_texture_module_n_177);
  vga_com_texture_module_g11276 : AO221D0BWP7T port map(A1 => vga_com_texture_module_n_140, A2 => vga_com_texture_module_n_15, B1 => vga_com_texture_module_n_144, B2 => vga_com_texture_module_hvis(2), C => vga_com_texture_module_n_168, Z => vga_com_texture_module_n_176);
  vga_com_texture_module_g11277 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_158, B1 => vga_com_column(0), B2 => FE_PHN17_vga_com_texture_module_n_20, ZN => vga_com_texture_module_n_175);
  vga_com_texture_module_g11278 : OAI222D0BWP7T port map(A1 => vga_com_texture_module_n_145, A2 => vga_com_texture_module_n_104, B1 => xplayer(1), B2 => vga_com_texture_module_n_120, C1 => vga_com_texture_module_n_102, C2 => vga_com_texture_module_n_141, ZN => vga_com_texture_module_n_174);
  vga_com_texture_module_g11279 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_128, B1 => vga_com_texture_module_n_167, ZN => vga_com_texture_module_n_182);
  vga_com_texture_module_g11280 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_167, A2 => vga_com_texture_module_n_128, ZN => vga_com_texture_module_n_180);
  vga_com_texture_module_g11281 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_156, A2 => vga_com_texture_module_n_84, A3 => FE_OFN0_reset, ZN => vga_com_texture_module_n_178);
  vga_com_texture_module_g11282 : HA1D0BWP7T port map(A => FE_PHN211_vga_com_hcount_6, B => vga_com_texture_module_n_133, CO => vga_com_texture_module_n_170, S => vga_com_texture_module_n_171);
  vga_com_texture_module_g11283 : INR2XD0BWP7T port map(A1 => vga_com_texture_module_n_158, B1 => vga_com_texture_module_n_142, ZN => vga_com_texture_module_n_173);
  vga_com_texture_module_g11284 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_158, A2 => vga_com_column(0), Z => vga_com_texture_module_n_172);
  vga_com_texture_module_g11292 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_140, A2 => vga_com_texture_module_n_77, B => vga_com_texture_module_n_155, Z => vga_com_texture_module_n_165);
  vga_com_texture_module_g11293 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_127, A2 => vga_com_texture_module_xposition(2), B1 => vga_com_texture_module_n_127, B2 => vga_com_texture_module_xposition(2), ZN => vga_com_texture_module_n_164);
  vga_com_texture_module_g11294 : IAO21D0BWP7T port map(A1 => vga_com_texture_module_n_145, A2 => vga_com_texture_module_n_76, B => vga_com_texture_module_n_160, ZN => vga_com_texture_module_n_163);
  vga_com_texture_module_g11295 : OAI31D0BWP7T port map(A1 => vga_com_texture_module_xposition(0), A2 => vga_com_texture_module_n_116, A3 => vga_com_texture_module_n_135, B => vga_com_texture_module_n_157, ZN => vga_com_texture_module_n_162);
  vga_com_texture_module_g11296 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_140, A2 => vga_com_texture_module_n_5, B1 => vga_com_texture_module_n_144, B2 => vga_com_texture_module_hvis(4), ZN => vga_com_texture_module_n_161);
  vga_com_texture_module_g11297 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_140, A2 => vga_com_texture_module_n_86, B1 => vga_com_texture_module_n_144, B2 => vga_com_texture_module_n_76, ZN => vga_com_texture_module_n_169);
  vga_com_texture_module_g11298 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_145, A2 => vga_com_texture_module_n_45, B1 => vga_com_texture_module_n_140, B2 => vga_com_texture_module_n_36, ZN => vga_com_texture_module_n_168);
  vga_com_texture_module_g11299 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_130, A2 => FE_OFN0_reset, B1 => vga_com_texture_module_n_143, B2 => vga_com_texture_module_n_108, ZN => vga_com_texture_module_n_167);
  vga_com_texture_module_g11300 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_156, B1 => FE_OFN0_reset, ZN => vga_com_texture_module_n_166);
  vga_com_texture_module_g11301 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_142, B1 => vga_com_texture_module_xposition(0), ZN => vga_com_texture_module_n_157);
  vga_com_texture_module_g11302 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_141, A2 => vga_com_texture_module_n_86, ZN => vga_com_texture_module_n_160);
  vga_com_texture_module_g11304 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_127, B1 => vga_com_texture_module_xposition(2), ZN => vga_com_texture_module_n_159);
  vga_com_texture_module_g11305 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_142, A2 => vga_com_texture_module_n_41, Z => vga_com_texture_module_n_158);
  vga_com_texture_module_g11307 : INVD1BWP7T port map(I => vga_com_texture_module_n_153, ZN => vga_com_texture_module_n_152);
  vga_com_texture_module_g11308 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_137, A2 => FE_OFN1_vga_com_row_0, B1 => vga_com_texture_module_n_137, B2 => FE_OFN1_vga_com_row_0, ZN => vga_com_texture_module_n_151);
  vga_com_texture_module_g11309 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_131, A2 => FE_PHN253_vga_com_texture_module_yposition_0, B1 => vga_com_texture_module_n_131, B2 => FE_PHN253_vga_com_texture_module_yposition_0, ZN => vga_com_texture_module_n_150);
  vga_com_texture_module_g11310 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_141, A2 => vga_com_texture_module_n_36, A3 => vga_com_texture_module_hvis(2), ZN => vga_com_texture_module_n_149);
  vga_com_texture_module_g11311 : IND4D0BWP7T port map(A1 => vga_com_texture_module_n_125, B1 => vga_com_hcount(5), B2 => FE_PHN235_vga_com_hcount_9, B3 => vga_com_texture_module_n_1, ZN => vga_com_texture_module_n_156);
  vga_com_texture_module_g11312 : AN3D0BWP7T port map(A1 => vga_com_texture_module_n_144, A2 => vga_com_texture_module_n_45, A3 => vga_com_texture_module_n_15, Z => vga_com_texture_module_n_155);
  vga_com_texture_module_g11313 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_135, A2 => vga_com_texture_module_n_91, B => vga_com_texture_module_n_84, ZN => vga_com_texture_module_n_154);
  vga_com_texture_module_g11314 : INR2D1BWP7T port map(A1 => vga_com_texture_module_n_108, B1 => vga_com_texture_module_n_143, ZN => vga_com_texture_module_n_153);
  vga_com_texture_module_g11315 : INVD1BWP7T port map(I => vga_com_texture_module_n_145, ZN => vga_com_texture_module_n_144);
  vga_com_texture_module_g11316 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_131, B1 => FE_PHN253_vga_com_texture_module_yposition_0, ZN => vga_com_texture_module_n_148);
  vga_com_texture_module_g11317 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_137, B1 => FE_OFN1_vga_com_row_0, ZN => vga_com_texture_module_n_147);
  vga_com_texture_module_g11318 : IOA21D1BWP7T port map(A1 => vga_com_texture_module_n_95, A2 => FE_DBTN0_reset, B => vga_com_texture_module_n_135, ZN => vga_com_texture_module_n_146);
  vga_com_texture_module_g11319 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_123, B1 => vga_com_texture_module_n_132, ZN => vga_com_texture_module_n_145);
  vga_com_texture_module_g11320 : INVD1BWP7T port map(I => vga_com_texture_module_n_141, ZN => vga_com_texture_module_n_140);
  vga_com_texture_module_g11321 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_114, A2 => vga_com_timer1(5), B1 => vga_com_texture_module_n_114, B2 => vga_com_timer1(5), ZN => vga_com_texture_module_n_138);
  vga_com_texture_module_g11322 : ND3D0BWP7T port map(A1 => vga_com_texture_module_n_126, A2 => vga_com_texture_module_n_37, A3 => FE_DBTN0_reset, ZN => vga_com_texture_module_n_143);
  vga_com_texture_module_g11323 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_136, A2 => vga_com_texture_module_n_116, ZN => vga_com_texture_module_n_142);
  vga_com_texture_module_g11324 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_132, A2 => vga_com_texture_module_n_123, ZN => vga_com_texture_module_n_141);
  vga_com_texture_module_g11325 : AOI31D1BWP7T port map(A1 => vga_com_texture_module_n_121, A2 => FE_PHN235_vga_com_hcount_9, A3 => vga_com_hcount(8), B => FE_OFN0_reset, ZN => vga_com_texture_module_n_139);
  vga_com_texture_module_g11326 : INVD1BWP7T port map(I => vga_com_texture_module_n_136, ZN => vga_com_texture_module_n_135);
  vga_com_texture_module_g11327 : HA1D0BWP7T port map(A => vga_com_hcount(5), B => vga_com_texture_module_n_117, CO => vga_com_texture_module_n_133, S => FE_PHN219_vga_com_texture_module_n_134);
  vga_com_texture_module_g11328 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_33, B1 => vga_com_texture_module_n_126, ZN => vga_com_texture_module_n_137);
  vga_com_texture_module_g11330 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_126, A2 => FE_OFN0_reset, ZN => vga_com_texture_module_n_136);
  vga_com_texture_module_g11331 : OAI211D1BWP7T port map(A1 => vga_com_texture_module_yposition(4), A2 => vga_com_texture_module_n_109, B => vga_com_texture_module_n_126, C => vga_com_texture_module_n_38, ZN => vga_com_texture_module_n_130);
  vga_com_texture_module_g11332 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_122, A2 => vga_com_texture_module_xposition(1), B1 => vga_com_texture_module_n_122, B2 => vga_com_texture_module_xposition(1), ZN => vga_com_texture_module_n_129);
  vga_com_texture_module_g11333 : NR2D1BWP7T port map(A1 => vga_com_texture_module_n_124, A2 => FE_OFN0_reset, ZN => vga_com_texture_module_n_132);
  vga_com_texture_module_g11334 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_85, B1 => vga_com_texture_module_n_126, ZN => vga_com_texture_module_n_131);
  vga_com_texture_module_g11335 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_26, A2 => FE_PHN239_vga_com_vcount_8, B => vga_com_texture_module_n_113, C => FE_PHN241_vga_com_vcount_9, ZN => vga_com_texture_module_n_128);
  vga_com_texture_module_g11336 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_122, B1 => vga_com_texture_module_xposition(1), ZN => vga_com_texture_module_n_127);
  vga_com_texture_module_g11337 : IND4D0BWP7T port map(A1 => vga_com_hcount(6), B1 => vga_com_hcount(4), B2 => vga_com_hcount(7), B3 => vga_com_texture_module_n_101, ZN => vga_com_texture_module_n_125);
  vga_com_texture_module_g11338 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_34, A2 => vga_com_texture_module_xposition(4), B => vga_com_texture_module_n_119, ZN => vga_com_texture_module_n_124);
  vga_com_texture_module_g11339 : AN4D1BWP7T port map(A1 => vga_com_texture_module_n_117, A2 => vga_com_texture_module_n_60, A3 => FE_PHN235_vga_com_hcount_9, A4 => vga_com_hcount(8), Z => vga_com_texture_module_n_126);
  vga_com_texture_module_g11340 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_116, A2 => vga_com_texture_module_n_60, ZN => vga_com_texture_module_n_121);
  vga_com_texture_module_g11341 : AOI211XD0BWP7T port map(A1 => vga_com_texture_module_n_98, A2 => vga_com_hcount(8), B => vga_com_texture_module_n_111, C => FE_PHN235_vga_com_hcount_9, ZN => vga_com_texture_module_n_123);
  vga_com_texture_module_g11342 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_117, A2 => vga_com_texture_module_xposition(0), ZN => vga_com_texture_module_n_122);
  vga_com_texture_module_g11343 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_80, A2 => vga_com_texture_module_n_67, B1 => vga_com_texture_module_n_112, B2 => vga_com_texture_module_n_34, ZN => vga_com_texture_module_n_119);
  vga_com_texture_module_g11344 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_97, A2 => vga_com_texture_module_timer1(4), B1 => vga_com_texture_module_n_97, B2 => vga_com_texture_module_timer1(4), ZN => vga_com_texture_module_n_118);
  vga_com_texture_module_g11345 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_34, B1 => FE_DBTN0_reset, B2 => vga_com_texture_module_n_112, ZN => vga_com_texture_module_n_120);
  vga_com_texture_module_g11346 : INVD1BWP7T port map(I => vga_com_texture_module_n_117, ZN => vga_com_texture_module_n_116);
  vga_com_texture_module_g11347 : HA1D0BWP7T port map(A => vga_com_hcount(4), B => vga_com_texture_module_n_99, CO => vga_com_texture_module_n_117, S => vga_com_texture_module_n_115);
  vga_com_texture_module_g11349 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_4, A2 => yplayer(3), B => vga_com_texture_module_n_110, ZN => vga_com_texture_module_n_113);
  vga_com_texture_module_g11350 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_97, B1 => vga_com_texture_module_timer1(4), ZN => vga_com_texture_module_n_114);
  vga_com_texture_module_g11351 : IAO21D0BWP7T port map(A1 => vga_com_texture_module_n_98, A2 => vga_com_hcount(8), B => xplayer(3), ZN => vga_com_texture_module_n_111);
  vga_com_texture_module_g11352 : INR4D0BWP7T port map(A1 => vga_com_texture_module_n_92, B1 => vga_com_hcount(8), B2 => vga_com_hcount(4), B3 => FE_PHN235_vga_com_hcount_9, ZN => vga_com_texture_module_n_112);
  vga_com_texture_module_g11353 : MAOI222D1BWP7T port map(A => vga_com_texture_module_n_87, B => vga_com_texture_module_n_27, C => vga_com_vcount(7), ZN => vga_com_texture_module_n_110);
  vga_com_texture_module_g11354 : OAI221D0BWP7T port map(A1 => vga_com_texture_module_n_7, A2 => yplayer(3), B1 => vga_com_texture_module_n_47, B2 => vga_com_texture_module_n_73, C => vga_com_texture_module_n_96, ZN => vga_com_texture_module_n_109);
  vga_com_texture_module_g11355 : INVD0BWP7T port map(I => vga_com_texture_module_n_106, ZN => vga_com_texture_module_n_107);
  vga_com_texture_module_g11356 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_74, A2 => vga_com_hcount(3), B => vga_com_texture_module_n_101, Z => FE_PHN197_vga_com_texture_module_n_105);
  vga_com_texture_module_g11357 : NR4D0BWP7T port map(A1 => vga_com_texture_module_n_83, A2 => FE_PHN241_vga_com_vcount_9, A3 => FE_PHN231_vga_com_vcount_2, A4 => vga_com_vcount(3), ZN => vga_com_texture_module_n_108);
  vga_com_texture_module_g11358 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_100, A2 => vga_com_texture_module_n_671, ZN => vga_com_texture_module_n_106);
  vga_com_texture_module_g11359 : XNR2D1BWP7T port map(A1 => vga_com_texture_module_n_89, A2 => vga_com_texture_module_hvis(6), ZN => vga_com_texture_module_n_104);
  vga_com_texture_module_g11360 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_72, A2 => vga_com_texture_module_timer1(3), B1 => vga_com_texture_module_n_72, B2 => vga_com_texture_module_timer1(3), ZN => vga_com_texture_module_n_103);
  vga_com_texture_module_g11361 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_93, A2 => vga_com_texture_module_hvis(6), B1 => vga_com_texture_module_n_93, B2 => vga_com_texture_module_hvis(6), ZN => vga_com_texture_module_n_102);
  vga_com_texture_module_g11362 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_74, A2 => vga_com_hcount(3), ZN => vga_com_texture_module_n_101);
  vga_com_texture_module_g11363 : INR2XD0BWP7T port map(A1 => vga_com_hcount(3), B1 => vga_com_texture_module_n_74, ZN => vga_com_texture_module_n_99);
  vga_com_texture_module_g11365 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_75, A2 => vga_com_texture_module_vvis(3), ZN => vga_com_texture_module_n_100);
  vga_com_texture_module_g11366 : AO31D1BWP7T port map(A1 => vga_com_texture_module_n_73, A2 => vga_com_texture_module_n_47, A3 => vga_com_texture_module_n_7, B => vga_com_texture_module_n_25, Z => vga_com_texture_module_n_96);
  vga_com_texture_module_g11367 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_83, B1 => FE_PHN241_vga_com_vcount_9, B2 => vga_com_texture_module_n_31, ZN => vga_com_texture_module_n_95);
  vga_com_texture_module_g11368 : OAI31D0BWP7T port map(A1 => xplayer(0), A2 => vga_com_texture_module_n_3, A3 => vga_com_texture_module_n_0, B => vga_com_texture_module_n_88, ZN => vga_com_texture_module_n_98);
  vga_com_texture_module_g11369 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_72, B1 => vga_com_texture_module_timer1(3), ZN => vga_com_texture_module_n_97);
  vga_com_texture_module_g11370 : INVD0BWP7T port map(I => vga_com_texture_module_n_75, ZN => vga_com_texture_module_n_94);
  vga_com_texture_module_g11371 : NR4D0BWP7T port map(A1 => vga_com_texture_module_n_66, A2 => vga_com_hcount(0), A3 => vga_com_hcount(3), A4 => vga_com_hcount(1), ZN => vga_com_texture_module_n_92);
  vga_com_texture_module_g11372 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_85, A2 => FE_DBTN0_reset, ZN => vga_com_texture_module_n_91);
  vga_com_texture_module_g11373 : OR2D1BWP7T port map(A1 => vga_com_texture_module_n_86, A2 => vga_com_texture_module_n_670, Z => vga_com_texture_module_n_93);
  vga_com_texture_module_g11374 : AOI222D0BWP7T port map(A1 => vga_com_texture_module_n_61, A2 => vga_com_hcount(4), B1 => vga_com_texture_module_n_24, B2 => vga_com_hcount(7), C1 => vga_com_texture_module_n_57, C2 => vga_com_hcount(6), ZN => vga_com_texture_module_n_88);
  vga_com_texture_module_g11375 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_78, A2 => vga_com_texture_module_vvis(5), A3 => vga_com_texture_module_vvis(4), ZN => vga_com_texture_module_n_90);
  vga_com_texture_module_g11376 : MAOI222D1BWP7T port map(A => vga_com_texture_module_n_64, B => yplayer(1), C => vga_com_texture_module_n_2, ZN => vga_com_texture_module_n_87);
  vga_com_texture_module_g11377 : NR3D0BWP7T port map(A1 => vga_com_texture_module_n_76, A2 => vga_com_texture_module_hvis(4), A3 => vga_com_texture_module_hvis(5), ZN => vga_com_texture_module_n_89);
  vga_com_texture_module_g11380 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_77, A2 => FE_PHN251_vga_com_texture_module_hvis_3, ZN => vga_com_texture_module_n_86);
  vga_com_texture_module_g11383 : IND3D1BWP7T port map(A1 => vga_com_texture_module_n_33, B1 => vga_com_vcount(4), B2 => vga_com_texture_module_n_31, ZN => vga_com_texture_module_n_85);
  vga_com_texture_module_g11384 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_35, A2 => vga_com_texture_module_timer1(2), B1 => vga_com_texture_module_n_35, B2 => vga_com_texture_module_timer1(2), ZN => vga_com_texture_module_n_82);
  vga_com_texture_module_g11385 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_44, A2 => vga_com_texture_module_vvis(2), B1 => vga_com_texture_module_n_44, B2 => vga_com_texture_module_vvis(2), ZN => vga_com_texture_module_n_81);
  vga_com_texture_module_g11386 : AOI221D0BWP7T port map(A1 => vga_com_texture_module_n_29, A2 => vga_com_texture_module_xposition(3), B1 => xplayer(2), B2 => vga_com_texture_module_xposition(2), C => vga_com_texture_module_n_65, ZN => vga_com_texture_module_n_80);
  vga_com_texture_module_g11387 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_n_41, A2 => vga_com_hcount(2), B1 => vga_com_texture_module_n_41, B2 => vga_com_hcount(2), ZN => vga_com_texture_module_n_79);
  vga_com_texture_module_g11388 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_63, A2 => vga_com_texture_module_n_32, B => vga_com_texture_module_n_19, ZN => vga_com_texture_module_n_84);
  vga_com_texture_module_g11389 : IND3D1BWP7T port map(A1 => vga_com_vcount(1), B1 => vga_com_texture_module_n_14, B2 => vga_com_texture_module_n_63, ZN => vga_com_texture_module_n_83);
  vga_com_texture_module_g11390 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_668, A2 => vga_com_texture_module_n_42, ZN => vga_com_texture_module_n_78);
  vga_com_texture_module_g11391 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_36, A2 => vga_com_texture_module_n_15, ZN => vga_com_texture_module_n_77);
  vga_com_texture_module_g11392 : ND2D1BWP7T port map(A1 => vga_com_texture_module_n_675, A2 => vga_com_texture_module_n_45, ZN => vga_com_texture_module_n_76);
  vga_com_texture_module_g11394 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_44, A2 => vga_com_texture_module_n_8, ZN => vga_com_texture_module_n_75);
  vga_com_texture_module_g11395 : IND2D1BWP7T port map(A1 => vga_com_texture_module_n_41, B1 => vga_com_hcount(2), ZN => vga_com_texture_module_n_74);
  vga_com_texture_module_g11396 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_58, A2 => vga_com_texture_module_frame_count(0), B => vga_com_texture_module_n_43, ZN => vga_com_texture_module_n_71);
  vga_com_texture_module_g11397 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_58, A2 => vga_com_texture_module_n_53, B => vga_com_texture_module_n_43, ZN => vga_com_texture_module_n_70);
  vga_com_texture_module_g11398 : IOA21D0BWP7T port map(A1 => vga_com_texture_module_n_59, A2 => vga_com_texture_module_n_682, B => vga_com_texture_module_n_43, ZN => vga_com_texture_module_n_69);
  vga_com_texture_module_g11399 : OAI22D0BWP7T port map(A1 => vga_com_texture_module_n_58, A2 => vga_com_texture_module_n_51, B1 => vga_com_texture_module_n_28, B2 => vga_com_texture_module_n_683, ZN => vga_com_texture_module_n_68);
  vga_com_texture_module_g11400 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_56, A2 => xplayer(3), B1 => vga_com_texture_module_n_24, B2 => xplayer(3), ZN => vga_com_texture_module_n_67);
  vga_com_texture_module_g11401 : OAI211D1BWP7T port map(A1 => vga_com_texture_module_yposition(2), A2 => yplayer(2), B => vga_com_texture_module_n_55, C => vga_com_texture_module_n_673, ZN => vga_com_texture_module_n_73);
  vga_com_texture_module_g11402 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_35, B1 => vga_com_texture_module_timer1(2), ZN => vga_com_texture_module_n_72);
  vga_com_texture_module_g11403 : IND2D1BWP7T port map(A1 => vga_com_hcount(2), B1 => vga_com_texture_module_n_60, ZN => vga_com_texture_module_n_66);
  vga_com_texture_module_g11404 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_672, A2 => vga_com_texture_module_n_30, B => vga_com_texture_module_n_669, ZN => vga_com_texture_module_n_65);
  vga_com_texture_module_g11405 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_40, A2 => yplayer(0), B => vga_com_texture_module_n_39, Z => vga_com_texture_module_n_64);
  vga_com_texture_module_g11406 : AOI32D1BWP7T port map(A1 => vga_com_texture_module_n_12, A2 => vga_com_column(1), A3 => vga_com_column(0), B1 => FE_PHN17_vga_com_texture_module_n_20, B2 => vga_com_column(2), ZN => vga_com_texture_module_n_62);
  vga_com_texture_module_g11407 : AOI21D0BWP7T port map(A1 => vga_com_texture_module_n_3, A2 => xplayer(0), B => vga_com_texture_module_n_0, ZN => vga_com_texture_module_n_61);
  vga_com_texture_module_g11408 : AN4D1BWP7T port map(A1 => vga_com_texture_module_n_39, A2 => vga_com_texture_module_n_10, A3 => vga_com_texture_module_n_2, A4 => vga_com_texture_module_n_4, Z => vga_com_texture_module_n_63);
  vga_com_texture_module_g11409 : CKND1BWP7T port map(I => vga_com_texture_module_n_58, ZN => vga_com_texture_module_n_59);
  vga_com_texture_module_g11410 : NR2D0BWP7T port map(A1 => vga_com_texture_module_n_46, A2 => xplayer(1), ZN => vga_com_texture_module_n_57);
  vga_com_texture_module_g11411 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_24, A2 => vga_com_texture_module_xposition(2), B => vga_com_texture_module_xposition(3), Z => vga_com_texture_module_n_56);
  vga_com_texture_module_g11412 : OAI21D0BWP7T port map(A1 => vga_com_texture_module_n_21, A2 => yplayer(0), B => vga_com_texture_module_n_674, ZN => vga_com_texture_module_n_55);
  vga_com_texture_module_g11414 : NR3D0BWP7T port map(A1 => vga_com_hcount(5), A2 => vga_com_hcount(6), A3 => vga_com_hcount(7), ZN => vga_com_texture_module_n_60);
  vga_com_texture_module_g11415 : AOI22D0BWP7T port map(A1 => vga_com_texture_module_n_678, A2 => vga_com_texture_module_n_681, B1 => vga_com_texture_module_n_679, B2 => vga_com_texture_module_n_683, ZN => vga_com_texture_module_n_58);
  vga_com_texture_module_g11416 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_712, A2 => vga_com_texture_module_frame_count(2), B1 => vga_com_texture_module_n_712, B2 => vga_com_texture_module_frame_count(2), ZN => vga_com_texture_module_n_53);
  vga_com_texture_module_g11417 : MOAI22D0BWP7T port map(A1 => FE_PHN199_vga_com_texture_module_n_18, A2 => vga_com_hcount(1), B1 => FE_PHN199_vga_com_texture_module_n_18, B2 => vga_com_hcount(1), ZN => vga_com_texture_module_n_52);
  vga_com_texture_module_g11418 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_676, A2 => vga_com_texture_module_frame_count(3), B1 => vga_com_texture_module_n_676, B2 => vga_com_texture_module_frame_count(3), ZN => vga_com_texture_module_n_51);
  vga_com_texture_module_g11419 : MAOI22D0BWP7T port map(A1 => yplayer(0), A2 => yplayer(1), B1 => yplayer(0), B2 => yplayer(1), ZN => vga_com_texture_module_n_50);
  vga_com_texture_module_g11420 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_14, A2 => vga_com_vcount(1), B1 => vga_com_texture_module_n_14, B2 => vga_com_vcount(1), ZN => vga_com_texture_module_n_49);
  vga_com_texture_module_g11421 : MAOI22D0BWP7T port map(A1 => vga_com_texture_module_n_16, A2 => vga_com_texture_module_vvis(1), B1 => vga_com_texture_module_n_16, B2 => vga_com_texture_module_vvis(1), ZN => vga_com_texture_module_n_54);
  vga_com_texture_module_g11422 : MAOI22D0BWP7T port map(A1 => FE_PHN193_vga_com_texture_module_n_17, A2 => vga_com_texture_module_hvis(1), B1 => FE_PHN193_vga_com_texture_module_n_17, B2 => vga_com_texture_module_hvis(1), ZN => vga_com_texture_module_n_48);
  vga_com_texture_module_g11424 : CKND2D1BWP7T port map(A1 => vga_com_vcount(4), A2 => vga_com_vcount(5), ZN => vga_com_texture_module_n_40);
  vga_com_texture_module_g11425 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_27, A2 => vga_com_texture_module_n_26, ZN => vga_com_texture_module_n_47);
  vga_com_texture_module_g11426 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_n_24, A2 => vga_com_hcount(7), ZN => vga_com_texture_module_n_46);
  vga_com_texture_module_g11427 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_hvis(0), A2 => vga_com_texture_module_hvis(1), ZN => vga_com_texture_module_n_45);
  vga_com_texture_module_g11428 : ND2D1BWP7T port map(A1 => vga_com_texture_module_vvis(1), A2 => vga_com_texture_module_vvis(0), ZN => vga_com_texture_module_n_44);
  vga_com_texture_module_g11429 : IND2D0BWP7T port map(A1 => vga_com_texture_module_n_681, B1 => vga_com_texture_module_n_678, ZN => vga_com_texture_module_n_43);
  vga_com_texture_module_g11430 : NR2XD0BWP7T port map(A1 => vga_com_texture_module_vvis(0), A2 => vga_com_texture_module_vvis(1), ZN => vga_com_texture_module_n_42);
  vga_com_texture_module_g11431 : ND2D1BWP7T port map(A1 => vga_com_hcount(0), A2 => vga_com_hcount(1), ZN => vga_com_texture_module_n_41);
  vga_com_texture_module_g11433 : INVD0BWP7T port map(I => vga_com_texture_module_n_37, ZN => vga_com_texture_module_n_38);
  vga_com_texture_module_g11434 : INVD0BWP7T port map(I => vga_com_texture_module_n_32, ZN => vga_com_texture_module_n_31);
  vga_com_texture_module_g11435 : IND2D0BWP7T port map(A1 => xplayer(0), B1 => vga_com_texture_module_xposition(0), ZN => vga_com_texture_module_n_30);
  vga_com_texture_module_g11436 : ND2D0BWP7T port map(A1 => xplayer(2), A2 => xplayer(3), ZN => vga_com_texture_module_n_29);
  vga_com_texture_module_g11437 : NR2XD0BWP7T port map(A1 => vga_com_vcount(4), A2 => vga_com_vcount(5), ZN => vga_com_texture_module_n_39);
  vga_com_texture_module_g11438 : NR2XD0BWP7T port map(A1 => yplayer(3), A2 => yplayer(2), ZN => vga_com_texture_module_n_37);
  vga_com_texture_module_g11439 : ND2D1BWP7T port map(A1 => vga_com_texture_module_hvis(1), A2 => vga_com_texture_module_hvis(0), ZN => vga_com_texture_module_n_36);
  vga_com_texture_module_g11440 : IND2D0BWP7T port map(A1 => vga_com_texture_module_timer1(1), B1 => vga_com_texture_module_timer1(0), ZN => vga_com_texture_module_n_35);
  vga_com_texture_module_g11441 : IND2D1BWP7T port map(A1 => xplayer(3), B1 => vga_com_texture_module_n_24, ZN => vga_com_texture_module_n_34);
  vga_com_texture_module_g11442 : ND2D1BWP7T port map(A1 => vga_com_vcount(1), A2 => vga_com_vcount(0), ZN => vga_com_texture_module_n_33);
  vga_com_texture_module_g11443 : ND2D1BWP7T port map(A1 => vga_com_vcount(3), A2 => FE_PHN231_vga_com_vcount_2, ZN => vga_com_texture_module_n_32);
  vga_com_texture_module_g11445 : INVD1BWP7T port map(I => yplayer(2), ZN => vga_com_texture_module_n_27);
  vga_com_texture_module_g11459 : INVD1BWP7T port map(I => yplayer(3), ZN => vga_com_texture_module_n_26);
  vga_com_texture_module_g11573 : INVD1BWP7T port map(I => xplayer(2), ZN => vga_com_texture_module_n_24);
  vga_com_texture_module_column_reg_1 : DFD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_206, Q => vga_com_column(1), QN => vga_com_texture_module_n_20);
  vga_com_texture_module_column_reg_2 : DFD1BWP7T port map(CP => CTS_23, D => FE_PHN298_vga_com_texture_module_n_202, Q => vga_com_column(2), QN => vga_com_texture_module_n_12);
  vga_com_texture_module_hcount_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN199_vga_com_texture_module_n_18, CP => CTS_23, D => vga_com_texture_module_n_139, Q => vga_com_hcount(0), QN => vga_com_texture_module_n_18);
  vga_com_texture_module_hcount_reg_5 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_134, CP => CTS_23, D => vga_com_texture_module_n_139, Q => vga_com_hcount(5), QN => vga_com_texture_module_n_3);
  vga_com_texture_module_hcount_reg_6 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_171, CP => CTS_23, D => vga_com_texture_module_n_139, Q => vga_com_hcount(6), QN => vga_com_texture_module_n_13);
  vga_com_texture_module_hcount_reg_8 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_139, CP => CTS_23, D => vga_com_texture_module_n_232, Q => FE_PHN236_vga_com_hcount_8, QN => vga_com_texture_module_n_1);
  vga_com_texture_module_hvis_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN193_vga_com_texture_module_n_17, CP => CTS_23, D => vga_com_texture_module_n_132, Q => vga_com_texture_module_hvis(0), QN => vga_com_texture_module_n_17);
  vga_com_texture_module_hvis_reg_2 : DFD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_216, Q => vga_com_texture_module_hvis(2), QN => vga_com_texture_module_n_15);
  vga_com_texture_module_hvis_reg_4 : DFD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_187, Q => vga_com_texture_module_hvis(4), QN => vga_com_texture_module_n_5);
  vga_com_texture_module_hvis_reg_5 : DFD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_223, Q => vga_com_texture_module_hvis(5), QN => vga_com_texture_module_n_22);
  vga_com_texture_module_timer1_reg_0 : DFCND1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_done, D => vga_com_texture_module_n_11, Q => vga_com_texture_module_timer1(0), QN => vga_com_texture_module_n_11);
  vga_com_texture_module_vcount_reg_0 : DFXD1BWP7T port map(CP => CTS_23, DA => vga_com_texture_module_n_166, DB => vga_com_texture_module_n_178, Q => vga_com_vcount(0), QN => vga_com_texture_module_n_14, SA => FE_PHN200_vga_com_vcount_0);
  vga_com_texture_module_vcount_reg_5 : DFD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_231, Q => FE_PHN242_vga_com_vcount_5, QN => vga_com_texture_module_n_6);
  vga_com_texture_module_vcount_reg_6 : DFXD1BWP7T port map(CP => CTS_23, DA => vga_com_texture_module_n_226, DB => vga_com_texture_module_n_192, Q => FE_PHN234_vga_com_vcount_6, QN => vga_com_texture_module_n_2, SA => vga_com_vcount(6));
  vga_com_texture_module_vcount_reg_7 : DFD1BWP7T port map(CP => CTS_23, D => FE_PHN281_vga_com_texture_module_n_244, Q => vga_com_vcount(7), QN => vga_com_texture_module_n_10);
  vga_com_texture_module_vcount_reg_8 : DFXD1BWP7T port map(CP => CTS_23, DA => vga_com_texture_module_n_235, DB => vga_com_texture_module_n_219, Q => vga_com_vcount(8), QN => vga_com_texture_module_n_4, SA => FE_PHN239_vga_com_vcount_8);
  vga_com_texture_module_vcount_reg_9 : DFD1BWP7T port map(CP => CTS_23, D => FE_PHN335_vga_com_texture_module_n_251, Q => vga_com_vcount(9), QN => vga_com_texture_module_n_19);
  vga_com_texture_module_vvis_reg_0 : DFD1BWP7T port map(CP => CTS_23, D => vga_com_texture_module_n_213, Q => FE_PHN252_vga_com_texture_module_vvis_0, QN => FE_PHN204_vga_com_texture_module_n_16);
  vga_com_texture_module_vvis_reg_2 : DFD1BWP7T port map(CP => CTS_23, D => FE_PHN339_vga_com_texture_module_n_249, Q => vga_com_texture_module_vvis(2), QN => vga_com_texture_module_n_8);
  vga_com_texture_module_vvis_reg_4 : DFD1BWP7T port map(CP => CTS_23, D => FE_PHN259_vga_com_texture_module_n_247, Q => vga_com_texture_module_vvis(4), QN => vga_com_texture_module_n_9);
  vga_com_texture_module_yposition_reg_0 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_150, CP => CTS_23, D => vga_com_texture_module_n_146, Q => vga_com_texture_module_yposition(0), QN => vga_com_texture_module_n_21);
  vga_com_texture_module_yposition_reg_2 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_146, CP => CTS_23, D => FE_PHN325_vga_com_texture_module_n_229, Q => vga_com_texture_module_yposition(2), QN => vga_com_texture_module_n_7);
  vga_com_texture_module_g2 : AO21D0BWP7T port map(A1 => vga_com_texture_module_n_13, A2 => xplayer(1), B => vga_com_texture_module_n_46, Z => vga_com_texture_module_n_0);
  vga_com_texture_module_g16998 : CKXOR2D1BWP7T port map(A1 => vga_com_texture_module_vvis(6), A2 => vga_com_texture_module_n_664, Z => vga_com_texture_module_n_850);
  vga_com_texture_module_timer1_reg_4 : DFCND1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_done, D => vga_com_texture_module_n_118, Q => vga_com_texture_module_timer1(4), QN => vga_com_texture_module_n_651);
  vga_com_texture_module_hvis_reg_1 : DFXD1BWP7T port map(CP => CTS_23, DA => vga_com_texture_module_n_144, DB => vga_com_texture_module_n_140, Q => vga_com_texture_module_hvis(1), QN => vga_com_texture_module_n_650, SA => FE_PHN326_vga_com_texture_module_n_48);
  vga_com_texture_module_yposition_reg_1 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_146, CP => CTS_23, D => FE_PHN361_vga_com_texture_module_n_190, Q => vga_com_texture_module_yposition(1), QN => vga_com_texture_module_n_266);
  vga_com_texture_module_xposition_reg_0 : DFD1BWP7T port map(CP => CTS_23, D => FE_PHN331_vga_com_texture_module_n_162, Q => vga_com_texture_module_xposition(0), QN => vga_com_texture_module_n_265);
  vga_com_texture_module_frame_count_reg_2 : DFCND1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_com_texture_module_timer1(4), D => vga_com_texture_module_n_70, Q => vga_com_texture_module_frame_count(2), QN => vga_com_texture_module_n_264);
  vga_com_texture_module_frame_count_reg_3 : DFCND1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_com_texture_module_timer1(4), D => vga_com_texture_module_n_68, Q => vga_com_texture_module_frame_count(3), QN => vga_com_texture_module_n_263);
  vga_com_texture_module_frame_count_reg_1 : DFCND1BWP7T port map(CDN => FE_DBTN0_reset, CP => vga_com_texture_module_timer1(4), D => vga_com_texture_module_n_69, Q => vga_com_texture_module_frame_count(1), QN => vga_com_texture_module_n_260);
  vga_com_texture_module_xposition_reg_2 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_136, CP => CTS_23, D => FE_PHN194_vga_com_texture_module_n_164, Q => vga_com_texture_module_xposition(2), QN => vga_com_texture_module_n_259);
  vga_com_texture_module_yposition_reg_3 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_146, CP => CTS_23, D => vga_com_texture_module_n_252, Q => vga_com_texture_module_yposition(3), QN => vga_com_texture_module_n_25);
  vga_com_texture_module_xposition_reg_3 : DFKCND1BWP7T port map(CN => vga_com_texture_module_n_136, CP => CTS_23, D => FE_PHN213_vga_com_texture_module_n_204, Q => vga_com_texture_module_xposition(3), QN => vga_com_texture_module_n_257);
  vga_com_texture_module_xposition_reg_1 : DFKCND1BWP7T port map(CN => FE_PHN386_vga_com_texture_module_n_129, CP => CTS_23, D => vga_com_texture_module_n_136, Q => vga_com_texture_module_xposition(1), QN => vga_com_texture_module_n_256);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1143 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_142, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_107, B1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_142, B2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_107, ZN => vga_com_texture_module_n_697);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1144 : MAOI222D1BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_140, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_115, C => vga_com_texture_module_csa_tree_add_99_11_groupi_n_96, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_142);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1145 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_140, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_118, B1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_140, B2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_118, ZN => vga_com_texture_module_n_696);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1146 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_125, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_114, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_137, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_140, S => vga_com_texture_module_n_695);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1147 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_126, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_127, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_135, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_137, S => vga_com_texture_module_n_694);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1148 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_128, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_121, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_133, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_135, S => vga_com_texture_module_n_693);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1149 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_122, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_119, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_131, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_133, S => vga_com_texture_module_n_692);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1150 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_120, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_108, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_129, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_131, S => vga_com_texture_module_n_691);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1151 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_109, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_101, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_123, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_129, S => vga_com_texture_module_n_690);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1152 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_112, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_89, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_111, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_127, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_128);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1153 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_110, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_91, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_104, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_125, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_126);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1154 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_116, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_84, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_102, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_123, S => vga_com_texture_module_n_689);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1155 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_105, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_90, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_113, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_121, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_122);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1156 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_64, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_97, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_106, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_119, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_120);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1157 : XNR2D1BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_115, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_96, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_118);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1158 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_99, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_70, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_85, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_116, S => vga_com_texture_module_n_688);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1159 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_77, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_71, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_103, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_115, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_114);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1160 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_93, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_63, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_83, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_112, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_113);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1161 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_68, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_82, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_92, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_110, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_111);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1162 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_62, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_74, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_98, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_108, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_109);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1163 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_95, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_59, B1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_95, B2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_59, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_107);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1164 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_73, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_61, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_94, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_105, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_106);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1165 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_57, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_67, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_72, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_103, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_104);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1166 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_54, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_69, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_81, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_101, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_102);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1167 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_50, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_65, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_86, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_99, S => vga_com_texture_module_n_687);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1168 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_53, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_52, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_80, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_97, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_98);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1169 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_79, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_78, B1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_79, B2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_78, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_96);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1170 : MAOI222D1BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_88, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_60, C => vga_com_texture_module_csa_tree_add_99_11_groupi_n_20, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_95);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1171 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_3, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_51, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_56, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_93, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_94);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1172 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_22, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_45, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_75, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_91, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_92);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1173 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_55, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_7, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_76, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_89, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_90);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1174 : INVD0BWP7T port map(I => vga_com_texture_module_csa_tree_add_99_11_groupi_n_78, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_88);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1175 : HA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_32, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_66, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_86, S => vga_com_texture_module_n_686);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1176 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_2, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_48, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_49, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_84, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_85);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1177 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_9, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_46, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_6, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_82, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_83);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1178 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_30, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_47, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_8, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_80, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_81);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1179 : CKXOR2D1BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_60, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_20, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_79);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1180 : MAOI222D1BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_58, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_40, C => vga_com_texture_module_csa_tree_add_99_11_groupi_n_41, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_78);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1181 : MOAI22D0BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_42, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_58, B1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_42, B2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_58, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_77);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1182 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_28, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_17, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_23, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_75, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_76);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1183 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_10, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_5, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_12, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_73, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_74);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1184 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_27, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_26, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_13, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_71, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_72);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1185 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_18, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_24, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_25, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_69, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_70);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1186 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_1, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_0, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_34, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_67, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_68);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1187 : FA1D0BWP7T port map(A => vga_com_texture_module_n_706, B => vga_com_texture_module_n_699, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_11, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_65, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_66);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1188 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_4, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_29, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_15, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_63, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_64);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1189 : FA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_21, B => vga_com_texture_module_n_708, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_36, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_61, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_62);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1190 : FA1D0BWP7T port map(A => vga_com_texture_module_n_850, B => vga_com_texture_module_n_711, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_37, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_59, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_60);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1191 : FA1D0BWP7T port map(A => vga_com_texture_module_n_710, B => vga_com_texture_module_n_703, CI => vga_com_texture_module_csa_tree_add_99_11_groupi_n_14, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_58, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_57);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1192 : HA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_38, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_31, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_55, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_56);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1193 : HA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_35, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_39, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_53, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_54);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1194 : HA1D0BWP7T port map(A => vga_com_texture_module_n_701, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_16, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_51, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_52);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1195 : HA1D0BWP7T port map(A => vga_com_texture_module_csa_tree_add_99_11_groupi_n_33, B => vga_com_texture_module_csa_tree_add_99_11_groupi_n_19, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_49, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_50);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1196 : HA1D0BWP7T port map(A => vga_com_texture_module_n_700, B => vga_com_texture_module_n_707, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_47, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_48);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1197 : HA1D0BWP7T port map(A => vga_com_texture_module_n_702, B => vga_com_texture_module_n_709, CO => vga_com_texture_module_csa_tree_add_99_11_groupi_n_45, S => vga_com_texture_module_csa_tree_add_99_11_groupi_n_46);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1198 : HA1D0BWP7T port map(A => vga_com_texture_module_n_705, B => vga_com_texture_module_n_698, CO => vga_com_texture_module_n_685, S => vga_com_texture_module_n_684);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1199 : XNR2D1BWP7T port map(A1 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_40, A2 => vga_com_texture_module_csa_tree_add_99_11_groupi_n_41, ZN => vga_com_texture_module_csa_tree_add_99_11_groupi_n_42);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1200 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_709, A2 => vga_com_texture_module_n_705, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_39);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1201 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_709, A2 => vga_com_texture_module_n_707, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_38);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1202 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_711, A2 => vga_com_texture_module_n_710, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_37);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1203 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_710, A2 => vga_com_texture_module_n_705, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_36);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1204 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_701, A2 => vga_com_texture_module_n_699, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_35);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1205 : AN2D0BWP7T port map(A1 => vga_com_texture_module_n_850, A2 => vga_com_texture_module_n_700, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_34);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1206 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_700, A2 => vga_com_texture_module_n_698, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_33);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1207 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_706, A2 => vga_com_texture_module_n_705, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_32);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1208 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_710, A2 => vga_com_texture_module_n_706, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_31);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1209 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_708, A2 => vga_com_texture_module_n_706, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_30);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1210 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_702, A2 => vga_com_texture_module_n_700, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_29);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1211 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_711, A2 => vga_com_texture_module_n_709, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_41);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1212 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_709, A2 => vga_com_texture_module_n_708, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_28);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1213 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_711, A2 => vga_com_texture_module_n_708, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_27);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1214 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_850, A2 => vga_com_texture_module_n_702, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_40);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1215 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_703, A2 => vga_com_texture_module_n_702, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_26);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1216 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_707, A2 => vga_com_texture_module_n_706, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_25);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1217 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_700, A2 => vga_com_texture_module_n_699, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_24);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1218 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_710, A2 => vga_com_texture_module_n_707, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_23);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1219 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_703, A2 => vga_com_texture_module_n_701, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_22);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1220 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_708, A2 => vga_com_texture_module_n_707, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_21);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1221 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_707, A2 => vga_com_texture_module_n_705, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_19);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1222 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_701, A2 => vga_com_texture_module_n_698, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_18);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1223 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_702, A2 => vga_com_texture_module_n_701, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_17);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1224 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_701, A2 => vga_com_texture_module_n_700, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_16);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1225 : AN2D0BWP7T port map(A1 => vga_com_texture_module_n_850, A2 => vga_com_texture_module_n_698, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_15);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1226 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_710, A2 => vga_com_texture_module_n_709, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_14);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1227 : AN2D0BWP7T port map(A1 => vga_com_texture_module_n_850, A2 => vga_com_texture_module_n_701, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_13);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1228 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_703, A2 => vga_com_texture_module_n_698, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_12);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1229 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_699, A2 => vga_com_texture_module_n_698, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_11);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1230 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_709, A2 => vga_com_texture_module_n_706, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_10);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1231 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_711, A2 => vga_com_texture_module_n_706, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_9);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1232 : AN2D0BWP7T port map(A1 => vga_com_texture_module_n_702, A2 => vga_com_texture_module_n_698, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_8);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1233 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_703, A2 => vga_com_texture_module_n_700, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_7);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1234 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_850, A2 => vga_com_texture_module_n_703, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_20);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1235 : AN2D0BWP7T port map(A1 => vga_com_texture_module_n_850, A2 => vga_com_texture_module_n_699, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_6);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1236 : AN2D1BWP7T port map(A1 => vga_com_texture_module_n_702, A2 => vga_com_texture_module_n_699, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_5);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1237 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_711, A2 => vga_com_texture_module_n_705, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_4);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1238 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_703, A2 => vga_com_texture_module_n_699, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_3);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1239 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_708, A2 => vga_com_texture_module_n_705, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_2);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1240 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_711, A2 => vga_com_texture_module_n_707, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_1);
  vga_com_texture_module_csa_tree_add_99_11_groupi_g1241 : CKAN2D1BWP7T port map(A1 => vga_com_texture_module_n_710, A2 => vga_com_texture_module_n_708, Z => vga_com_texture_module_csa_tree_add_99_11_groupi_n_0);
  vga_com_tile_module_g47695 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_93, A2 => vga_com_tile_module_n_1015, B => vga_com_tile_module_n_1041, C => vga_com_tile_module_n_988, ZN => vga_com_color_address(0));
  vga_com_tile_module_g47696 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_1040, A2 => vga_com_tile_module_n_99, B1 => vga_com_tile_module_n_1014, B2 => vga_com_tile_module_n_240, ZN => vga_com_tile_module_n_1041);
  vga_com_tile_module_g47697 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_1039, A2 => vga_com_tile_address(4), B1 => vga_com_tile_module_n_98, B2 => vga_com_tile_module_n_1007, C1 => vga_com_tile_module_n_96, C2 => vga_com_tile_module_n_985, ZN => vga_com_tile_module_n_1040);
  vga_com_tile_module_g47698 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_6, A2 => vga_com_tile_module_n_869, A3 => vga_com_tile_module_n_54, B => vga_com_tile_module_n_1038, ZN => vga_com_tile_module_n_1039);
  vga_com_tile_module_g47699 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_1033, A2 => vga_com_tile_module_n_6, B1 => vga_com_tile_module_n_963, B2 => vga_com_tile_module_n_89, ZN => vga_com_tile_module_n_1038);
  vga_com_tile_module_g47700 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_1034, A2 => vga_com_tile_module_n_93, B1 => vga_com_tile_module_n_1023, B2 => vga_com_tile_module_n_99, ZN => vga_com_color_address(3));
  vga_com_tile_module_g47701 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_1031, A2 => vga_com_tile_module_n_93, B1 => vga_com_tile_module_n_1009, B2 => vga_com_tile_module_n_99, ZN => vga_com_color_address(2));
  vga_com_tile_module_g47702 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_1027, A2 => vga_com_tile_address(5), B => vga_com_tile_module_n_1022, C => FE_OFN0_reset, Z => vga_com_color_address(1));
  vga_com_tile_module_g47703 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_55, A2 => vga_com_tile_module_n_747, A3 => vga_com_tile_module_n_94, B => vga_com_tile_module_n_1030, ZN => vga_com_tile_module_n_1034);
  vga_com_tile_module_g47704 : OAI32D1BWP7T port map(A1 => vga_com_tile_module_n_998, A2 => vga_com_tile_module_n_858, A3 => vga_com_tile_module_n_49, B1 => vga_com_tile_address(2), B2 => vga_com_tile_module_n_1028, ZN => vga_com_tile_module_n_1033);
  vga_com_tile_module_g47705 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_93, A2 => vga_com_tile_module_n_97, A3 => vga_com_tile_module_n_996, B => vga_com_tile_module_n_1029, ZN => vga_com_color_address(4));
  vga_com_tile_module_g47706 : OA221D0BWP7T port map(A1 => vga_com_tile_module_n_1024, A2 => vga_com_tile_address(4), B1 => vga_com_tile_module_n_98, B2 => vga_com_tile_module_n_968, C => vga_com_tile_module_n_1018, Z => vga_com_tile_module_n_1031);
  vga_com_tile_module_g47707 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_97, A2 => vga_com_tile_module_n_1003, B => vga_com_tile_module_n_1025, C => vga_com_tile_module_n_758, ZN => vga_com_tile_module_n_1030);
  vga_com_tile_module_g47708 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_994, A2 => vga_com_tile_module_n_99, B1 => vga_com_tile_module_n_1026, B2 => vga_com_tile_module_n_93, ZN => vga_com_tile_module_n_1029);
  vga_com_tile_module_g47709 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_1021, A2 => vga_com_tile_module_n_3, B1 => vga_com_tile_module_n_992, B2 => vga_com_tile_address(1), C => vga_com_tile_module_n_402, ZN => vga_com_tile_module_n_1028);
  vga_com_tile_module_g47710 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_976, A2 => vga_com_tile_module_n_98, B1 => vga_com_tile_module_n_97, B2 => vga_com_tile_module_n_983, C => vga_com_tile_module_n_1016, ZN => vga_com_tile_module_n_1027);
  vga_com_tile_module_g47711 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_1020, A2 => vga_com_tile_address(4), B1 => vga_com_tile_module_n_990, B2 => vga_com_tile_module_n_94, ZN => vga_com_tile_module_n_1026);
  vga_com_tile_module_g47712 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_1017, A2 => vga_com_tile_address(4), B1 => vga_com_tile_module_n_924, B2 => vga_com_tile_module_n_214, ZN => vga_com_tile_module_n_1025);
  vga_com_tile_module_g47713 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_1000, A2 => vga_com_tile_module_n_6, B => vga_com_tile_module_n_949, C => vga_com_tile_module_n_941, ZN => vga_com_tile_module_n_1024);
  vga_com_tile_module_g47714 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_68, A2 => vga_com_tile_module_n_995, B => vga_com_tile_module_n_1019, C => vga_com_tile_module_n_1008, ZN => vga_com_tile_module_n_1023);
  vga_com_tile_module_g47715 : AN3D0BWP7T port map(A1 => vga_com_tile_module_n_1013, A2 => vga_com_tile_module_n_83, A3 => vga_com_tile_module_n_94, Z => vga_com_tile_module_n_1022);
  vga_com_tile_module_g47716 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_124, A2 => vga_com_tile_module_n_182, B => vga_com_tile_module_n_1011, C => vga_com_tile_module_n_533, ZN => vga_com_tile_module_n_1021);
  vga_com_tile_module_g47717 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_993, A2 => vga_com_tile_address(3), B1 => vga_com_tile_module_n_842, B2 => vga_com_tile_module_n_241, C => vga_com_tile_module_n_999, ZN => vga_com_tile_module_n_1020);
  vga_com_tile_module_g47718 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_425, A2 => vga_com_tile_module_n_68, B => vga_com_tile_module_n_1005, C => vga_com_tile_module_n_230, ZN => vga_com_tile_module_n_1019);
  vga_com_tile_module_g47719 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_981, A2 => vga_com_tile_module_n_89, A3 => vga_com_tile_address(4), B => vga_com_tile_module_n_1012, ZN => vga_com_tile_module_n_1018);
  vga_com_tile_module_g47720 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_1002, A2 => vga_com_tile_address(3), B1 => vga_com_tile_module_n_95, B2 => vga_com_tile_module_n_982, C1 => vga_com_tile_module_n_90, C2 => vga_com_tile_module_n_971, ZN => vga_com_tile_module_n_1017);
  vga_com_tile_module_g47721 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_970, A2 => vga_com_tile_module_n_94, B1 => vga_com_tile_module_n_1004, B2 => vga_com_tile_module_n_96, ZN => vga_com_tile_module_n_1016);
  vga_com_tile_module_g47722 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_1001, A2 => vga_com_tile_module_n_13, B => vga_com_tile_module_n_1010, ZN => vga_com_tile_module_n_1015);
  vga_com_tile_module_g47723 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_1006, A2 => vga_com_tile_address(2), B1 => vga_com_tile_module_n_86, B2 => vga_com_tile_module_n_904, ZN => vga_com_tile_module_n_1014);
  vga_com_tile_module_g47724 : NR4D0BWP7T port map(A1 => vga_com_tile_module_n_946, A2 => vga_com_tile_module_n_920, A3 => vga_com_tile_module_n_980, A4 => vga_com_tile_address(5), ZN => vga_com_tile_module_n_1013);
  vga_com_tile_module_g47725 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_979, A2 => vga_com_tile_module_n_917, A3 => vga_com_tile_module_n_987, B => vga_com_tile_module_n_96, ZN => vga_com_tile_module_n_1012);
  vga_com_tile_module_g47726 : ND3D0BWP7T port map(A1 => vga_com_tile_module_n_997, A2 => vga_com_tile_module_n_587, A3 => vga_com_tile_module_n_804, ZN => vga_com_tile_module_n_1011);
  vga_com_tile_module_g47727 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_984, A2 => vga_com_tile_module_n_870, B => vga_com_tile_module_n_96, ZN => vga_com_tile_module_n_1010);
  vga_com_tile_module_g47728 : OAI33D1BWP7T port map(A1 => vga_com_tile_module_n_229, A2 => vga_com_tile_module_n_967, A3 => vga_com_tile_module_n_977, B1 => vga_com_tile_module_n_959, B2 => vga_com_tile_address(1), B3 => vga_com_tile_module_n_214, ZN => vga_com_tile_module_n_1009);
  vga_com_tile_module_g47729 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_616, A2 => vga_com_tile_module_n_285, B => vga_com_tile_module_n_995, C => vga_com_tile_address(1), Z => vga_com_tile_module_n_1008);
  vga_com_tile_module_g47730 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_49, A2 => vga_com_tile_module_n_938, B => vga_com_tile_module_n_989, C => vga_com_tile_module_n_882, ZN => vga_com_tile_module_n_1007);
  vga_com_tile_module_g47731 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_906, A2 => vga_com_tile_module_n_60, B => vga_com_tile_module_n_885, C => vga_com_tile_module_n_978, ZN => vga_com_tile_module_n_1006);
  vga_com_tile_module_g47732 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_955, A2 => vga_com_tile_module_n_3, B1 => vga_com_tile_module_n_956, B2 => vga_com_tile_module_n_45, C => vga_com_tile_module_n_920, ZN => vga_com_tile_module_n_1005);
  vga_com_tile_module_g47733 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_45, A2 => vga_com_tile_address(2), A3 => vga_com_tile_module_n_573, B => vga_com_tile_module_n_986, ZN => vga_com_tile_module_n_1004);
  vga_com_tile_module_g47734 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_227, A2 => vga_com_tile_module_n_853, B => vga_com_tile_module_n_991, ZN => vga_com_tile_module_n_1003);
  vga_com_tile_module_g47735 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_950, A2 => vga_com_tile_address(2), B1 => vga_com_tile_module_n_86, B2 => vga_com_tile_module_n_907, C1 => vga_com_tile_module_n_952, C2 => vga_com_tile_module_n_55, ZN => vga_com_tile_module_n_1002);
  vga_com_tile_module_g47736 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_964, A2 => vga_com_tile_address(3), B1 => vga_com_tile_module_n_90, B2 => vga_com_tile_module_n_916, C1 => vga_com_tile_module_n_95, C2 => vga_com_tile_module_n_878, ZN => vga_com_tile_module_n_1001);
  vga_com_tile_module_g47737 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_49, A2 => vga_com_tile_module_n_925, B1 => vga_com_tile_module_n_975, B2 => vga_com_tile_module_n_83, C1 => vga_com_tile_module_n_854, C2 => vga_com_tile_module_n_54, ZN => vga_com_tile_module_n_1000);
  vga_com_tile_module_g47738 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_974, A2 => vga_com_tile_module_n_89, B1 => vga_com_tile_module_n_812, B2 => vga_com_tile_module_n_95, ZN => vga_com_tile_module_n_999);
  vga_com_tile_module_g47739 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_969, A2 => FE_OFN2_vga_com_tile_address_0, B1 => vga_com_tile_module_n_718, B2 => vga_com_tile_module_n_343, ZN => vga_com_tile_module_n_998);
  vga_com_tile_module_g47740 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_958, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_139, B2 => vga_com_tile_module_n_264, C1 => vga_com_tile_module_n_351, C2 => vga_com_tile_module_n_79, ZN => vga_com_tile_module_n_997);
  vga_com_tile_module_g47741 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_237, A2 => vga_com_tile_module_n_636, B1 => vga_com_tile_module_n_55, B2 => vga_com_tile_module_n_619, C => vga_com_tile_module_n_965, ZN => vga_com_tile_module_n_996);
  vga_com_tile_module_g47742 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_214, A2 => vga_com_tile_module_n_934, B => vga_com_tile_module_n_910, C => vga_com_tile_module_n_915, ZN => vga_com_tile_module_n_994);
  vga_com_tile_module_g47743 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_942, A2 => vga_com_tile_module_n_5, B => vga_com_tile_module_n_933, C => vga_com_tile_module_n_880, ZN => vga_com_tile_module_n_993);
  vga_com_tile_module_g47744 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_943, A2 => FE_OFN2_vga_com_tile_address_0, B => vga_com_tile_module_n_750, C => vga_com_tile_module_n_864, ZN => vga_com_tile_module_n_992);
  vga_com_tile_module_g47745 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_745, A2 => vga_com_tile_module_n_83, B => vga_com_tile_module_n_947, C => vga_com_tile_module_n_795, ZN => vga_com_tile_module_n_991);
  vga_com_tile_module_g47746 : AO222D0BWP7T port map(A1 => vga_com_tile_module_n_953, A2 => vga_com_tile_address(2), B1 => vga_com_tile_module_n_237, B2 => vga_com_tile_module_n_827, C1 => vga_com_tile_module_n_785, C2 => vga_com_tile_module_n_86, Z => vga_com_tile_module_n_990);
  vga_com_tile_module_g47747 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_898, A2 => vga_com_tile_module_n_37, B => vga_com_tile_module_n_973, ZN => vga_com_tile_module_n_995);
  vga_com_tile_module_g47748 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_954, A2 => vga_com_tile_module_n_5, B1 => vga_com_tile_module_n_158, B2 => vga_com_tile_module_n_752, ZN => vga_com_tile_module_n_989);
  vga_com_tile_module_g47749 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_951, A2 => vga_com_tile_module_n_417, B => vga_com_tile_module_n_54, C => vga_com_tile_module_n_240, Z => vga_com_tile_module_n_988);
  vga_com_tile_module_g47750 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_48, A2 => vga_com_tile_module_n_921, A3 => vga_com_tile_module_n_189, A4 => vga_com_tile_module_n_136, ZN => vga_com_tile_module_n_987);
  vga_com_tile_module_g47751 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_33, A2 => vga_com_tile_module_n_760, A3 => vga_com_tile_module_n_49, B => vga_com_tile_module_n_972, ZN => vga_com_tile_module_n_986);
  vga_com_tile_module_g47752 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_848, A2 => vga_com_tile_module_n_49, B => vga_com_tile_module_n_769, C => vga_com_tile_module_n_966, ZN => vga_com_tile_module_n_985);
  vga_com_tile_module_g47753 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_957, A2 => vga_com_tile_address(2), B1 => vga_com_tile_module_n_902, B2 => vga_com_tile_module_n_86, C1 => vga_com_tile_module_n_55, C2 => vga_com_tile_module_n_908, ZN => vga_com_tile_module_n_984);
  vga_com_tile_module_g47754 : AOI32D1BWP7T port map(A1 => vga_com_tile_module_n_863, A2 => vga_com_tile_module_n_859, A3 => vga_com_tile_module_n_5, B1 => vga_com_tile_module_n_962, B2 => vga_com_tile_address(2), ZN => vga_com_tile_module_n_983);
  vga_com_tile_module_g47755 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_918, A2 => vga_com_tile_address(1), B => vga_com_tile_module_n_834, C => vga_com_tile_module_n_903, ZN => vga_com_tile_module_n_982);
  vga_com_tile_module_g47756 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_236, A2 => vga_com_tile_module_n_896, B1 => vga_com_tile_module_n_764, B2 => vga_com_tile_address(1), C => vga_com_tile_module_n_948, ZN => vga_com_tile_module_n_981);
  vga_com_tile_module_g47757 : AOI221D0BWP7T port map(A1 => FE_PDN7_vga_com_tile_module_n_914, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_698, B2 => FE_OFN2_vga_com_tile_address_0, C => vga_com_tile_module_n_5, ZN => vga_com_tile_module_n_980);
  vga_com_tile_module_g47758 : OAI211D1BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_909, B => vga_com_tile_module_n_765, C => vga_com_tile_module_n_5, ZN => vga_com_tile_module_n_979);
  vga_com_tile_module_g47759 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_2, A2 => vga_com_tile_module_n_936, B => vga_com_tile_address(1), ZN => vga_com_tile_module_n_978);
  vga_com_tile_module_g47760 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_935, A2 => vga_com_tile_address(1), A3 => vga_com_tile_module_n_456, ZN => vga_com_tile_module_n_977);
  vga_com_tile_module_g47761 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_227, A2 => vga_com_tile_module_n_702, A3 => vga_com_tile_module_n_16, B => vga_com_tile_module_n_961, ZN => vga_com_tile_module_n_976);
  vga_com_tile_module_g47762 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_191, A2 => vga_com_tile_module_n_180, A3 => vga_com_tile_module_n_136, B => vga_com_tile_module_n_960, ZN => vga_com_tile_module_n_975);
  vga_com_tile_module_g47763 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_803, A2 => vga_com_tile_module_n_42, B => vga_com_tile_module_n_890, C => vga_com_tile_module_n_940, ZN => vga_com_tile_module_n_974);
  vga_com_tile_module_g47764 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_919, A2 => vga_com_tile_module_n_749, A3 => vga_com_tile_module_n_39, B => vga_com_tile_module_n_214, ZN => vga_com_tile_module_n_973);
  vga_com_tile_module_g47765 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_881, A2 => vga_com_tile_address(1), B => vga_com_tile_module_n_928, C => vga_com_tile_module_n_5, ZN => vga_com_tile_module_n_972);
  vga_com_tile_module_g47766 : AOI22D0BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_923, B1 => vga_com_tile_module_n_69, B2 => vga_com_tile_module_n_873, ZN => vga_com_tile_module_n_971);
  vga_com_tile_module_g47767 : NR4D0BWP7T port map(A1 => vga_com_tile_module_n_766, A2 => vga_com_tile_module_n_705, A3 => vga_com_tile_module_n_868, A4 => vga_com_tile_module_n_932, ZN => vga_com_tile_module_n_970);
  vga_com_tile_module_g47768 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_893, A2 => vga_com_tile_module_n_9, B => vga_com_tile_module_n_750, C => vga_com_tile_module_n_284, ZN => vga_com_tile_module_n_969);
  vga_com_tile_module_g47769 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_86, A2 => vga_com_tile_module_n_875, B1 => vga_com_tile_module_n_55, B2 => vga_com_tile_module_n_931, ZN => vga_com_tile_module_n_968);
  vga_com_tile_module_g47770 : OAI32D1BWP7T port map(A1 => vga_com_tile_module_n_174, A2 => vga_com_tile_module_n_44, A3 => vga_com_tile_module_n_905, B1 => vga_com_tile_module_n_820, B2 => vga_com_tile_module_n_70, ZN => vga_com_tile_module_n_967);
  vga_com_tile_module_g47771 : AOI32D1BWP7T port map(A1 => vga_com_tile_module_n_912, A2 => vga_com_tile_module_n_877, A3 => vga_com_tile_module_n_5, B1 => vga_com_tile_module_n_82, B2 => vga_com_tile_module_n_825, ZN => vga_com_tile_module_n_966);
  vga_com_tile_module_g47772 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_666, A2 => vga_com_tile_module_n_83, B => vga_com_tile_module_n_937, C => vga_com_tile_module_n_788, ZN => vga_com_tile_module_n_965);
  vga_com_tile_module_g47773 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_922, A2 => vga_com_tile_module_n_5, B1 => vga_com_tile_address(2), B2 => vga_com_tile_module_n_888, C1 => vga_com_tile_module_n_899, C2 => vga_com_tile_module_n_242, ZN => vga_com_tile_module_n_964);
  vga_com_tile_module_g47774 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_44, A2 => vga_com_tile_module_n_663, B => vga_com_tile_module_n_929, ZN => vga_com_tile_module_n_963);
  vga_com_tile_module_g47775 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_268, A2 => vga_com_tile_module_n_42, B => vga_com_tile_module_n_891, C => vga_com_tile_module_n_665, ZN => vga_com_tile_module_n_962);
  vga_com_tile_module_g47776 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_792, A2 => vga_com_tile_address(2), A3 => vga_com_tile_module_n_68, B => vga_com_tile_module_n_926, ZN => vga_com_tile_module_n_961);
  vga_com_tile_module_g47777 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_627, A2 => vga_com_tile_module_n_34, B1 => vga_com_tile_module_n_124, B2 => vga_com_tile_module_n_198, C => vga_com_tile_module_n_944, ZN => vga_com_tile_module_n_960);
  vga_com_tile_module_g47778 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_778, A2 => vga_com_tile_module_n_37, B1 => vga_com_tile_module_n_2, B2 => vga_com_tile_module_n_724, C => vga_com_tile_module_n_930, ZN => vga_com_tile_module_n_959);
  vga_com_tile_module_g47779 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_669, A2 => vga_com_tile_module_n_110, B1 => vga_com_tile_module_n_470, B2 => vga_com_tile_module_n_568, C => vga_com_tile_module_n_939, ZN => vga_com_tile_module_n_958);
  vga_com_tile_module_g47780 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_71, A2 => vga_com_tile_module_n_170, B => vga_com_tile_module_n_927, C => vga_com_tile_module_n_845, ZN => vga_com_tile_module_n_957);
  vga_com_tile_module_g47781 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_886, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_tile_module_n_299, B2 => vga_com_tile_module_n_633, C1 => vga_com_tile_module_n_18, C2 => vga_com_tile_module_n_577, ZN => vga_com_tile_module_n_956);
  vga_com_tile_module_g47782 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_887, A2 => vga_com_tile_module_n_33, B => vga_com_tile_module_n_686, C => vga_com_tile_module_n_456, Z => vga_com_tile_module_n_955);
  vga_com_tile_module_g47783 : OAI222D0BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_879, B1 => vga_com_tile_module_n_800, B2 => vga_com_tile_module_n_70, C1 => vga_com_tile_module_n_851, C2 => vga_com_tile_module_n_44, ZN => vga_com_tile_module_n_954);
  vga_com_tile_module_g47784 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_43, A2 => vga_com_tile_module_n_646, B => vga_com_tile_module_n_824, C => vga_com_tile_module_n_895, ZN => vga_com_tile_module_n_953);
  vga_com_tile_module_g47785 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_871, A2 => vga_com_tile_module_n_499, A3 => vga_com_tile_module_n_406, A4 => vga_com_tile_module_n_354, ZN => vga_com_tile_module_n_952);
  vga_com_tile_module_g47786 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_282, A2 => vga_com_tile_module_n_259, B1 => vga_com_tile_module_n_292, B2 => vga_com_tile_module_n_338, C => vga_com_tile_module_n_911, ZN => vga_com_tile_module_n_951);
  vga_com_tile_module_g47787 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_913, A2 => vga_com_tile_module_n_3, B1 => vga_com_tile_module_n_838, B2 => vga_com_tile_module_n_797, ZN => vga_com_tile_module_n_950);
  vga_com_tile_module_g47788 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_901, A2 => vga_com_tile_module_n_90, B1 => vga_com_tile_module_n_814, B2 => vga_com_tile_module_n_95, ZN => vga_com_tile_module_n_949);
  vga_com_tile_module_g47789 : AOI33D1BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_33, A3 => vga_com_tile_module_n_865, B1 => vga_com_tile_module_n_69, B2 => vga_com_tile_module_n_259, B3 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_948);
  vga_com_tile_module_g47790 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_900, A2 => vga_com_tile_module_n_5, B1 => vga_com_tile_module_n_86, B2 => vga_com_tile_module_n_731, ZN => vga_com_tile_module_n_947);
  vga_com_tile_module_g47791 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_856, A2 => vga_com_tile_module_n_817, A3 => vga_com_tile_module_n_3, B => vga_com_tile_module_n_945, ZN => vga_com_tile_module_n_946);
  vga_com_tile_module_g47792 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_808, A2 => vga_com_tile_module_n_19, B1 => vga_com_tile_module_n_268, B2 => vga_com_tile_module_n_688, C => vga_com_tile_module_n_86, ZN => vga_com_tile_module_n_945);
  vga_com_tile_module_g47793 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_143, A2 => vga_com_tile_module_n_328, B1 => vga_com_tile_module_n_337, B2 => vga_com_tile_module_n_107, C => vga_com_tile_module_n_897, ZN => vga_com_tile_module_n_944);
  vga_com_tile_module_g47794 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_884, A2 => FE_OFN4_vga_com_row_2, B => vga_com_tile_module_n_285, ZN => vga_com_tile_module_n_943);
  vga_com_tile_module_g47795 : OAI32D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_833, A3 => vga_com_tile_module_n_844, B1 => vga_com_tile_module_n_2, B2 => vga_com_tile_module_n_866, ZN => vga_com_tile_module_n_942);
  vga_com_tile_module_g47796 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_839, A2 => vga_com_tile_module_n_645, A3 => vga_com_tile_module_n_372, B => vga_com_tile_module_n_241, ZN => vga_com_tile_module_n_941);
  vga_com_tile_module_g47797 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_805, A2 => vga_com_tile_module_n_528, B => vga_com_tile_module_n_71, C => vga_com_tile_module_n_0, ZN => vga_com_tile_module_n_940);
  vga_com_tile_module_g47798 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_658, A2 => vga_com_tile_module_n_295, B1 => vga_com_tile_module_n_675, B2 => vga_com_tile_module_n_17, C => vga_com_tile_module_n_892, ZN => vga_com_tile_module_n_939);
  vga_com_tile_module_g47799 : NR4D0BWP7T port map(A1 => vga_com_tile_module_n_835, A2 => vga_com_tile_module_n_593, A3 => vga_com_tile_module_n_131, A4 => vga_com_tile_module_n_137, ZN => vga_com_tile_module_n_938);
  vga_com_tile_module_g47800 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_872, A2 => vga_com_tile_module_n_45, B => vga_com_tile_address(2), ZN => vga_com_tile_module_n_937);
  vga_com_tile_module_g47801 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_661, A2 => vga_com_tile_module_n_301, A3 => vga_com_tile_module_n_815, B => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_936);
  vga_com_tile_module_g47802 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_122, A2 => vga_com_tile_module_n_852, B => vga_com_tile_module_n_773, C => vga_com_tile_module_n_534, ZN => vga_com_tile_module_n_935);
  vga_com_tile_module_g47803 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_3, A2 => vga_com_tile_module_n_719, A3 => vga_com_tile_module_n_0, B => vga_com_tile_module_n_889, ZN => vga_com_tile_module_n_934);
  vga_com_tile_module_g47804 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_867, A2 => vga_com_tile_module_n_480, A3 => vga_com_tile_module_n_807, B => vga_com_tile_module_n_49, ZN => vga_com_tile_module_n_933);
  vga_com_tile_module_g47805 : AOI31D0BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_816, A3 => vga_com_tile_module_n_678, B => vga_com_tile_address(2), ZN => vga_com_tile_module_n_932);
  vga_com_tile_module_g47806 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_108, A2 => vga_com_tile_module_n_171, B => vga_com_tile_module_n_860, C => vga_com_tile_module_n_672, ZN => vga_com_tile_module_n_931);
  vga_com_tile_module_g47807 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_852, A2 => vga_com_tile_module_n_2, A3 => vga_com_tile_module_n_28, B => vga_com_tile_module_n_821, ZN => vga_com_tile_module_n_930);
  vga_com_tile_module_g47808 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_71, A2 => vga_com_tile_module_n_840, B1 => vga_com_tile_module_n_3, B2 => vga_com_tile_module_n_806, C1 => vga_com_tile_module_n_69, C2 => vga_com_tile_module_n_802, ZN => vga_com_tile_module_n_929);
  vga_com_tile_module_g47809 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_453, A2 => vga_com_tile_module_n_108, A3 => vga_com_tile_module_n_823, B => vga_com_tile_address(1), ZN => vga_com_tile_module_n_928);
  vga_com_tile_module_g47810 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_876, A2 => vga_com_tile_address(1), B1 => vga_com_tile_module_n_60, B2 => vga_com_tile_module_n_754, ZN => vga_com_tile_module_n_927);
  vga_com_tile_module_g47811 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_158, A2 => vga_com_tile_module_n_883, B1 => vga_com_tile_module_n_242, B2 => vga_com_tile_module_n_692, ZN => vga_com_tile_module_n_926);
  vga_com_tile_module_g47812 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_32, A2 => vga_com_tile_module_n_410, A3 => vga_com_tile_module_n_520, B => vga_com_tile_module_n_894, ZN => vga_com_tile_module_n_925);
  vga_com_tile_module_g47813 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_69, A2 => vga_com_tile_module_n_747, B1 => vga_com_tile_module_n_45, B2 => vga_com_tile_module_n_715, C => vga_com_tile_module_n_874, ZN => vga_com_tile_module_n_924);
  vga_com_tile_module_g47814 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_709, A2 => vga_com_tile_module_n_189, B1 => vga_com_tile_module_n_830, B2 => vga_com_tile_module_n_32, C1 => vga_com_tile_module_n_796, C2 => vga_com_tile_module_n_107, ZN => vga_com_tile_module_n_923);
  vga_com_tile_module_g47815 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_69, A2 => vga_com_tile_module_n_829, B1 => vga_com_tile_module_n_43, B2 => vga_com_tile_module_n_846, C1 => vga_com_tile_module_n_855, C2 => vga_com_tile_address(1), ZN => vga_com_tile_module_n_922);
  vga_com_tile_module_g47816 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_33, A2 => vga_com_tile_module_n_179, B1 => vga_com_tile_module_n_810, B2 => vga_com_tile_module_n_2, C1 => vga_com_tile_module_n_34, C2 => vga_com_tile_module_n_329, ZN => vga_com_tile_module_n_921);
  vga_com_tile_module_g47817 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_755, A2 => vga_com_tile_module_n_156, A3 => vga_com_tile_module_n_10, B => vga_com_tile_module_n_732, ZN => vga_com_tile_module_n_919);
  vga_com_tile_module_g47818 : OAI211D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_791, B => vga_com_tile_module_n_708, C => vga_com_tile_module_n_417, ZN => vga_com_tile_module_n_918);
  vga_com_tile_module_g47819 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_82, A2 => vga_com_tile_module_n_787, A3 => vga_com_tile_module_n_2, A4 => vga_com_tile_module_n_110, ZN => vga_com_tile_module_n_917);
  vga_com_tile_module_g47820 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_43, A2 => vga_com_tile_module_n_567, B => vga_com_tile_module_n_822, C => vga_com_tile_module_n_813, ZN => vga_com_tile_module_n_916);
  vga_com_tile_module_g47821 : IND3D1BWP7T port map(A1 => vga_com_tile_module_n_97, B1 => vga_com_tile_module_n_826, B2 => vga_com_tile_module_n_86, ZN => vga_com_tile_module_n_915);
  vga_com_tile_module_g47822 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_720, A2 => vga_com_tile_module_n_9, B1 => vga_com_tile_module_n_268, B2 => vga_com_tile_module_n_772, C1 => vga_com_tile_module_n_464, C2 => vga_com_tile_module_n_474, ZN => vga_com_tile_module_n_914);
  vga_com_tile_module_g47823 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_283, A2 => vga_com_tile_module_n_34, B => vga_com_tile_module_n_849, C => vga_com_tile_module_n_753, ZN => vga_com_tile_module_n_913);
  vga_com_tile_module_g47824 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_637, A2 => FE_OFN2_vga_com_tile_address_0, B1 => vga_com_tile_module_n_2, B2 => vga_com_tile_module_n_782, C => vga_com_tile_module_n_3, ZN => vga_com_tile_module_n_912);
  vga_com_tile_module_g47825 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_368, A2 => vga_com_tile_module_n_335, B1 => vga_com_tile_module_n_65, B2 => vga_com_tile_module_n_129, C => vga_com_tile_module_n_861, ZN => vga_com_tile_module_n_911);
  vga_com_tile_module_g47826 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_771, A2 => vga_com_tile_module_n_69, B => vga_com_tile_module_n_230, C => vga_com_tile_module_n_0, ZN => vga_com_tile_module_n_910);
  vga_com_tile_module_g47827 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_121, A2 => vga_com_tile_module_n_169, B => vga_com_tile_module_n_847, C => vga_com_tile_module_n_478, ZN => vga_com_tile_module_n_909);
  vga_com_tile_module_g47828 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_153, A2 => vga_com_tile_module_n_290, B1 => vga_com_tile_module_n_358, B2 => vga_com_tile_module_n_134, C => vga_com_tile_module_n_857, ZN => vga_com_tile_module_n_908);
  vga_com_tile_module_g47829 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_518, A2 => vga_com_tile_module_n_819, A3 => vga_com_tile_module_n_513, A4 => vga_com_tile_module_n_157, ZN => vga_com_tile_module_n_907);
  vga_com_tile_module_g47830 : OA221D0BWP7T port map(A1 => vga_com_tile_module_n_21, A2 => vga_com_tile_module_n_574, B1 => vga_com_tile_module_n_24, B2 => vga_com_tile_module_n_259, C => vga_com_tile_module_n_862, Z => vga_com_tile_module_n_906);
  vga_com_tile_module_g47831 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_557, A2 => vga_com_tile_module_n_427, B => vga_com_tile_module_n_832, C => vga_com_tile_module_n_682, ZN => vga_com_tile_module_n_905);
  vga_com_tile_module_g47832 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_789, A2 => vga_com_tile_module_n_105, A3 => vga_com_tile_module_n_104, B => vga_com_tile_module_n_70, ZN => vga_com_tile_module_n_920);
  vga_com_tile_module_g47833 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_37, A2 => vga_com_tile_module_n_547, B => vga_com_tile_module_n_836, C => vga_com_tile_module_n_536, ZN => vga_com_tile_module_n_904);
  vga_com_tile_module_g47834 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_757, A2 => vga_com_tile_module_n_507, A3 => vga_com_tile_module_n_16, B => vga_com_tile_module_n_68, ZN => vga_com_tile_module_n_903);
  vga_com_tile_module_g47835 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_32, A2 => vga_com_tile_module_n_776, B => vga_com_tile_module_n_843, C => vga_com_tile_module_n_620, ZN => vga_com_tile_module_n_902);
  vga_com_tile_module_g47836 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_69, A2 => vga_com_tile_module_n_841, B1 => vga_com_tile_module_n_43, B2 => vga_com_tile_module_n_654, C1 => vga_com_tile_module_n_71, C2 => vga_com_tile_module_n_624, ZN => vga_com_tile_module_n_901);
  vga_com_tile_module_g47837 : AO222D0BWP7T port map(A1 => vga_com_tile_module_n_45, A2 => vga_com_tile_module_n_798, B1 => vga_com_tile_module_n_71, B2 => vga_com_tile_module_n_715, C1 => vga_com_tile_module_n_799, C2 => vga_com_tile_module_n_43, Z => vga_com_tile_module_n_900);
  vga_com_tile_module_g47838 : AOI221D1BWP7T port map(A1 => vga_com_tile_module_n_259, A2 => vga_com_tile_module_n_103, B1 => vga_com_tile_module_n_212, B2 => vga_com_tile_module_n_28, C => vga_com_tile_module_n_831, ZN => vga_com_tile_module_n_899);
  vga_com_tile_module_g47839 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_424, A2 => vga_com_tile_module_n_179, B1 => vga_com_tile_module_n_24, B2 => vga_com_tile_module_n_314, C => vga_com_tile_module_n_809, ZN => vga_com_tile_module_n_898);
  vga_com_tile_module_g47840 : OA222D0BWP7T port map(A1 => vga_com_tile_module_n_761, A2 => FE_OFN2_vga_com_tile_address_0, B1 => vga_com_tile_module_n_67, B2 => vga_com_tile_module_n_150, C1 => vga_com_tile_module_n_263, C2 => vga_com_tile_module_n_354, Z => vga_com_tile_module_n_897);
  vga_com_tile_module_g47841 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_426, A2 => vga_com_tile_module_n_781, B1 => vga_com_tile_module_n_578, B2 => vga_com_tile_module_n_181, C1 => vga_com_tile_module_n_338, C2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_896);
  vga_com_tile_module_g47842 : OAI32D1BWP7T port map(A1 => vga_com_tile_module_n_178, A2 => vga_com_tile_module_n_169, A3 => vga_com_tile_module_n_3, B1 => vga_com_tile_module_n_827, B2 => vga_com_tile_module_n_68, ZN => vga_com_tile_module_n_895);
  vga_com_tile_module_g47843 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_854, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_644, B2 => vga_com_tile_module_n_34, ZN => vga_com_tile_module_n_894);
  vga_com_tile_module_g47844 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_850, A2 => vga_com_tile_module_n_10, B1 => vga_com_tile_module_n_21, B2 => vga_com_tile_module_n_669, C => vga_com_tile_module_n_770, ZN => vga_com_tile_module_n_893);
  vga_com_tile_module_g47845 : OAI32D1BWP7T port map(A1 => vga_com_tile_module_n_118, A2 => vga_com_tile_module_n_183, A3 => vga_com_tile_module_n_270, B1 => vga_com_tile_module_n_29, B2 => vga_com_tile_module_n_850, ZN => vga_com_tile_module_n_892);
  vga_com_tile_module_g47846 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_69, A2 => vga_com_tile_module_n_853, B1 => vga_com_tile_module_n_71, B2 => vga_com_tile_module_n_746, ZN => vga_com_tile_module_n_891);
  vga_com_tile_module_g47847 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_45, A2 => vga_com_tile_module_n_828, B1 => vga_com_tile_module_n_69, B2 => vga_com_tile_module_n_748, ZN => vga_com_tile_module_n_890);
  vga_com_tile_module_g47848 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_44, A2 => vga_com_tile_module_n_800, B1 => vga_com_tile_module_n_70, B2 => vga_com_tile_module_n_851, ZN => vga_com_tile_module_n_889);
  vga_com_tile_module_g47849 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_71, A2 => vga_com_tile_module_n_829, B1 => vga_com_tile_module_n_69, B2 => vga_com_tile_module_n_828, ZN => vga_com_tile_module_n_888);
  vga_com_tile_module_g47850 : INVD0BWP7T port map(I => vga_com_tile_module_n_886, ZN => vga_com_tile_module_n_887);
  vga_com_tile_module_g47851 : OAI31D0BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_352, A3 => vga_com_tile_module_n_697, B => vga_com_tile_module_n_3, ZN => vga_com_tile_module_n_885);
  vga_com_tile_module_g47852 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_735, A2 => vga_com_tile_module_n_273, B1 => vga_com_tile_module_n_794, B2 => vga_com_tile_module_n_712, ZN => vga_com_tile_module_n_884);
  vga_com_tile_module_g47853 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_267, A2 => vga_com_tile_module_n_779, B => vga_com_tile_module_n_573, Z => vga_com_tile_module_n_883);
  vga_com_tile_module_g47854 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_131, A2 => vga_com_tile_module_n_615, A3 => vga_com_tile_module_n_736, B => vga_com_tile_module_n_82, ZN => vga_com_tile_module_n_882);
  vga_com_tile_module_g47855 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_413, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_160, B2 => vga_com_tile_module_n_73, C => vga_com_tile_module_n_818, ZN => vga_com_tile_module_n_881);
  vga_com_tile_module_g47856 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_683, A2 => vga_com_tile_module_n_484, A3 => vga_com_tile_module_n_797, B => vga_com_tile_module_n_83, ZN => vga_com_tile_module_n_880);
  vga_com_tile_module_g47857 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_837, A2 => vga_com_tile_module_n_291, ZN => vga_com_tile_module_n_879);
  vga_com_tile_module_g47858 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_68, A2 => vga_com_tile_module_n_70, B => vga_com_tile_module_n_855, Z => vga_com_tile_module_n_878);
  vga_com_tile_module_g47859 : IND4D0BWP7T port map(A1 => vga_com_tile_module_n_137, B1 => vga_com_tile_module_n_130, B2 => vga_com_tile_module_n_707, B3 => vga_com_tile_address(1), ZN => vga_com_tile_module_n_877);
  vga_com_tile_module_g47860 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_524, A2 => vga_com_tile_module_n_33, B => vga_com_tile_module_n_763, C => vga_com_tile_module_n_756, ZN => vga_com_tile_module_n_876);
  vga_com_tile_module_g47861 : NR4D0BWP7T port map(A1 => vga_com_tile_module_n_790, A2 => vga_com_tile_module_n_691, A3 => vga_com_tile_module_n_303, A4 => vga_com_tile_module_n_492, ZN => vga_com_tile_module_n_875);
  vga_com_tile_module_g47862 : OAI33D0BWP7T port map(A1 => vga_com_tile_module_n_370, A2 => vga_com_tile_module_n_740, A3 => vga_com_tile_module_n_42, B1 => vga_com_tile_module_n_63, B2 => vga_com_tile_module_n_20, B3 => vga_com_tile_module_n_236, ZN => vga_com_tile_module_n_874);
  vga_com_tile_module_g47863 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_706, A2 => vga_com_tile_module_n_594, A3 => vga_com_tile_module_n_459, A4 => vga_com_tile_module_n_247, ZN => vga_com_tile_module_n_873);
  vga_com_tile_module_g47864 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_564, A2 => vga_com_tile_address(1), B => vga_com_tile_module_n_759, C => vga_com_tile_module_n_665, ZN => vga_com_tile_module_n_872);
  vga_com_tile_module_g47865 : OAI211D1BWP7T port map(A1 => FE_OFN3_vga_com_row_1, A2 => vga_com_tile_module_n_727, B => vga_com_tile_module_n_749, C => vga_com_tile_module_n_703, ZN => vga_com_tile_module_n_886);
  vga_com_tile_module_g47866 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_137, A2 => vga_com_tile_module_n_190, B => vga_com_tile_module_n_385, C => vga_com_tile_module_n_767, ZN => vga_com_tile_module_n_871);
  vga_com_tile_module_g47867 : OAI31D1BWP7T port map(A1 => vga_com_tile_module_n_352, A2 => vga_com_tile_module_n_711, A3 => vga_com_tile_module_n_679, B => vga_com_tile_module_n_237, ZN => vga_com_tile_module_n_870);
  vga_com_tile_module_g47868 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_320, A2 => vga_com_tile_module_n_9, B => vga_com_tile_module_n_801, C => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_869);
  vga_com_tile_module_g47869 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_695, A2 => vga_com_tile_module_n_126, A3 => vga_com_tile_module_n_678, B => vga_com_tile_module_n_49, ZN => vga_com_tile_module_n_868);
  vga_com_tile_module_g47870 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_131, A2 => vga_com_column(1), B1 => vga_com_tile_module_n_733, B2 => vga_com_tile_module_n_34, C1 => vga_com_tile_module_n_135, C2 => vga_com_tile_module_n_85, ZN => vga_com_tile_module_n_867);
  vga_com_tile_module_g47871 : OAI33D1BWP7T port map(A1 => vga_com_tile_module_n_629, A2 => vga_com_tile_module_n_716, A3 => vga_com_tile_address(1), B1 => vga_com_tile_module_n_640, B2 => vga_com_tile_module_n_662, B3 => vga_com_tile_module_n_3, ZN => vga_com_tile_module_n_866);
  vga_com_tile_module_g47872 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_427, A2 => vga_com_tile_module_n_690, B1 => vga_com_tile_module_n_10, B2 => vga_com_tile_module_n_428, C1 => vga_com_tile_module_n_261, C2 => vga_com_tile_module_n_248, ZN => vga_com_tile_module_n_865);
  vga_com_tile_module_g47873 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_793, A2 => vga_com_tile_module_n_209, B1 => vga_com_tile_module_n_568, B2 => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_864);
  vga_com_tile_module_g47874 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_69, A2 => vga_com_tile_module_n_559, B1 => vga_com_tile_module_n_42, B2 => vga_com_tile_module_n_799, ZN => vga_com_tile_module_n_863);
  vga_com_tile_module_g47875 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_704, A2 => vga_com_tile_module_n_22, B1 => vga_com_tile_module_n_660, B2 => vga_com_tile_module_n_91, C1 => vga_com_tile_module_n_132, C2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_862);
  vga_com_tile_module_g47876 : OA221D0BWP7T port map(A1 => vga_com_tile_module_n_738, A2 => FE_OFN2_vga_com_tile_address_0, B1 => vga_com_tile_module_n_157, B2 => vga_com_tile_module_n_418, C => vga_com_tile_module_n_386, Z => vga_com_tile_module_n_861);
  vga_com_tile_module_g47877 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_189, A2 => vga_com_tile_module_n_333, B1 => vga_com_tile_module_n_37, B2 => vga_com_tile_module_n_693, C1 => vga_com_tile_module_n_2, C2 => vga_com_tile_module_n_550, ZN => vga_com_tile_module_n_860);
  vga_com_tile_module_g47878 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_71, A2 => vga_com_tile_module_n_580, B1 => vga_com_tile_module_n_44, B2 => vga_com_tile_module_n_798, ZN => vga_com_tile_module_n_859);
  vga_com_tile_module_g47879 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_278, A2 => vga_com_tile_module_n_125, B => vga_com_tile_module_n_741, C => vga_com_tile_module_n_768, ZN => vga_com_tile_module_n_858);
  vga_com_tile_module_g47880 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_676, A2 => vga_com_tile_module_n_203, B1 => vga_com_tile_module_n_776, B2 => vga_com_tile_module_n_38, ZN => vga_com_tile_module_n_857);
  vga_com_tile_module_g47881 : OA31D1BWP7T port map(A1 => vga_com_tile_module_n_41, A2 => vga_com_tile_module_n_196, A3 => vga_com_tile_module_n_153, B => vga_com_tile_module_n_811, Z => vga_com_tile_module_n_856);
  vga_com_tile_module_g47882 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_721, A2 => vga_com_tile_module_n_597, A3 => vga_com_tile_module_n_486, A4 => vga_com_tile_module_n_157, ZN => vga_com_tile_module_n_849);
  vga_com_tile_module_g47883 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_673, A2 => vga_com_tile_module_n_33, B => vga_com_tile_module_n_775, ZN => vga_com_tile_module_n_848);
  vga_com_tile_module_g47884 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_728, A2 => FE_OFN2_vga_com_tile_address_0, B => vga_com_tile_module_n_608, C => vga_com_tile_module_n_479, ZN => vga_com_tile_module_n_847);
  vga_com_tile_module_g47885 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_780, A2 => vga_com_tile_module_n_110, ZN => vga_com_tile_module_n_846);
  vga_com_tile_module_g47886 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_3, A2 => vga_com_tile_module_n_734, A3 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_845);
  vga_com_tile_module_g47887 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_611, A2 => vga_com_tile_module_n_9, B => vga_com_tile_address(1), C => vga_com_tile_module_n_542, ZN => vga_com_tile_module_n_844);
  vga_com_tile_module_g47888 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_676, A2 => vga_com_tile_module_n_108, B => vga_com_tile_module_n_783, C => vga_com_tile_module_n_556, ZN => vga_com_tile_module_n_843);
  vga_com_tile_module_g47889 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_108, A2 => vga_com_tile_module_n_319, B => vga_com_tile_module_n_672, C => vga_com_tile_module_n_680, ZN => vga_com_tile_module_n_842);
  vga_com_tile_module_g47890 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_466, A2 => vga_com_tile_module_n_18, B1 => vga_com_tile_module_n_26, B2 => vga_com_tile_module_n_363, C => vga_com_tile_module_n_777, ZN => vga_com_tile_module_n_841);
  vga_com_tile_module_g47891 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_670, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_tile_module_n_437, B2 => vga_com_tile_module_n_444, C => vga_com_tile_module_n_434, ZN => vga_com_tile_module_n_840);
  vga_com_tile_module_g47892 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_641, A2 => vga_com_tile_module_n_39, B1 => vga_com_tile_module_n_128, B2 => vga_com_tile_module_n_79, C => vga_com_tile_module_n_613, ZN => vga_com_tile_module_n_839);
  vga_com_tile_module_g47893 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_17, A2 => vga_com_tile_module_n_648, A3 => vga_com_tile_module_n_3, B => vga_com_tile_module_n_70, ZN => vga_com_tile_module_n_838);
  vga_com_tile_module_g47894 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_222, A2 => vga_com_tile_module_n_435, B => vga_com_tile_module_n_713, C => vga_com_tile_module_n_774, ZN => vga_com_tile_module_n_837);
  vga_com_tile_module_g47895 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_744, A2 => vga_com_tile_module_n_39, B => vga_com_tile_module_n_700, ZN => vga_com_tile_module_n_836);
  vga_com_tile_module_g47896 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_1, A2 => vga_com_tile_module_n_38, B1 => vga_com_tile_module_n_443, B2 => vga_com_tile_module_n_122, C => vga_com_tile_module_n_726, ZN => vga_com_tile_module_n_835);
  vga_com_tile_module_g47897 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_684, A2 => vga_com_tile_module_n_575, B => vga_com_tile_module_n_42, ZN => vga_com_tile_module_n_834);
  vga_com_tile_module_g47898 : NR4D0BWP7T port map(A1 => vga_com_tile_module_n_3, A2 => vga_com_tile_module_n_662, A3 => vga_com_tile_module_n_629, A4 => vga_com_tile_module_n_384, ZN => vga_com_tile_module_n_833);
  vga_com_tile_module_g47899 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_751, A2 => vga_com_tile_module_n_315, B => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_832);
  vga_com_tile_module_g47900 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_16, A2 => vga_com_tile_module_n_144, A3 => vga_com_tile_module_n_132, B => vga_com_tile_module_n_786, ZN => vga_com_tile_module_n_831);
  vga_com_tile_module_g47901 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_25, A2 => vga_com_tile_module_n_88, B => vga_com_tile_module_n_554, C => vga_com_tile_module_n_762, ZN => vga_com_tile_module_n_830);
  vga_com_tile_module_g47902 : ND3D0BWP7T port map(A1 => vga_com_tile_module_n_737, A2 => vga_com_tile_module_n_369, A3 => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_855);
  vga_com_tile_module_g47903 : AOI221D1BWP7T port map(A1 => vga_com_tile_module_n_664, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_tile_module_n_346, B2 => vga_com_tile_module_n_111, C => vga_com_tile_module_n_722, ZN => vga_com_tile_module_n_854);
  vga_com_tile_module_g47904 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_112, A2 => vga_com_tile_module_n_314, B => vga_com_tile_module_n_777, C => vga_com_tile_module_n_531, ZN => vga_com_tile_module_n_853);
  vga_com_tile_module_g47905 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_565, A2 => FE_OFN1_vga_com_row_0, B => vga_com_tile_module_n_751, C => vga_com_tile_module_n_199, ZN => vga_com_tile_module_n_852);
  vga_com_tile_module_g47906 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_395, A2 => vga_com_tile_module_n_320, B => vga_com_tile_module_n_801, ZN => vga_com_tile_module_n_851);
  vga_com_tile_module_g47907 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_743, A2 => FE_OFN1_vga_com_row_0, B => vga_com_tile_module_n_784, ZN => vga_com_tile_module_n_850);
  vga_com_tile_module_g47908 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_538, A2 => vga_com_tile_module_n_23, B1 => vga_com_tile_module_n_670, B2 => vga_com_tile_module_n_39, C1 => vga_com_tile_module_n_663, C2 => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_826);
  vga_com_tile_module_g47909 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_38, A2 => vga_com_tile_module_n_674, B => vga_com_tile_module_n_713, C => vga_com_tile_module_n_642, ZN => vga_com_tile_module_n_825);
  vga_com_tile_module_g47910 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_44, A2 => vga_com_tile_module_n_739, B1 => vga_com_tile_module_n_70, B2 => vga_com_tile_module_n_647, ZN => vga_com_tile_module_n_824);
  vga_com_tile_module_g47911 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_746, A2 => FE_OFN2_vga_com_tile_address_0, B1 => vga_com_tile_module_n_319, B2 => vga_com_tile_module_n_35, ZN => vga_com_tile_module_n_823);
  vga_com_tile_module_g47912 : OAI22D0BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_699, B1 => vga_com_tile_module_n_60, B2 => vga_com_tile_module_n_694, ZN => vga_com_tile_module_n_822);
  vga_com_tile_module_g47913 : AOI211D0BWP7T port map(A1 => vga_com_tile_module_n_62, A2 => vga_com_tile_module_n_50, B => vga_com_tile_module_n_689, C => vga_com_tile_module_n_152, ZN => vga_com_tile_module_n_821);
  vga_com_tile_module_g47914 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_630, A2 => vga_com_tile_module_n_523, A3 => vga_com_tile_module_n_105, A4 => vga_com_tile_module_n_114, ZN => vga_com_tile_module_n_820);
  vga_com_tile_module_g47915 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_160, A2 => vga_com_tile_module_n_223, B => vga_com_tile_module_n_305, C => vga_com_tile_module_n_701, ZN => vga_com_tile_module_n_819);
  vga_com_tile_module_g47916 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_746, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_183, B2 => vga_com_tile_module_n_162, ZN => vga_com_tile_module_n_818);
  vga_com_tile_module_g47917 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_725, A2 => vga_com_tile_module_n_370, B => vga_com_tile_module_n_267, Z => vga_com_tile_module_n_817);
  vga_com_tile_module_g47918 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_730, A2 => vga_com_tile_module_n_34, B1 => vga_com_tile_module_n_609, B2 => vga_com_tile_module_n_33, ZN => vga_com_tile_module_n_816);
  vga_com_tile_module_g47919 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_22, A2 => vga_com_tile_module_n_657, B1 => vga_com_tile_module_n_660, B2 => vga_com_tile_module_n_319, C1 => vga_com_tile_module_n_658, C2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_815);
  vga_com_tile_module_g47920 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_43, A2 => vga_com_tile_module_n_717, B1 => vga_com_tile_module_n_69, B2 => vga_com_tile_module_n_723, ZN => vga_com_tile_module_n_814);
  vga_com_tile_module_g47921 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_521, A2 => vga_com_tile_module_n_677, A3 => FE_OFN2_vga_com_tile_address_0, B => vga_com_tile_module_n_3, ZN => vga_com_tile_module_n_813);
  vga_com_tile_module_g47922 : AOI32D1BWP7T port map(A1 => vga_com_tile_module_n_69, A2 => vga_com_tile_module_n_656, A3 => vga_com_tile_module_n_63, B1 => vga_com_tile_module_n_43, B2 => vga_com_tile_module_n_639, ZN => vga_com_tile_module_n_812);
  vga_com_tile_module_g47923 : OA222D0BWP7T port map(A1 => vga_com_tile_module_n_149, A2 => vga_com_tile_module_n_337, B1 => vga_com_tile_module_n_37, B2 => vga_com_tile_module_n_671, C1 => vga_com_tile_module_n_38, C2 => vga_com_tile_module_n_650, Z => vga_com_tile_module_n_811);
  vga_com_tile_module_g47924 : AOI222D1BWP7T port map(A1 => vga_com_tile_module_n_634, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_tile_module_n_225, B2 => vga_com_tile_module_n_28, C1 => vga_com_tile_module_n_266, C2 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_810);
  vga_com_tile_module_g47925 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_667, A2 => vga_com_tile_module_n_20, B1 => vga_com_tile_module_n_571, B2 => vga_com_tile_module_n_22, C1 => vga_com_tile_module_n_356, C2 => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_809);
  vga_com_tile_module_g47926 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_268, A2 => vga_com_tile_module_n_2, B => vga_com_tile_module_n_729, C => vga_com_tile_module_n_283, Z => vga_com_tile_module_n_808);
  vga_com_tile_module_g47927 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_685, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_472, B2 => vga_com_tile_module_n_123, ZN => vga_com_tile_module_n_807);
  vga_com_tile_module_g47928 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_714, A2 => vga_com_tile_module_n_35, B1 => vga_com_tile_module_n_1, B2 => vga_com_tile_module_n_32, ZN => vga_com_tile_module_n_806);
  vga_com_tile_module_g47929 : OAI22D1BWP7T port map(A1 => vga_com_tile_module_n_16, A2 => vga_com_tile_module_n_668, B1 => vga_com_tile_module_n_18, B2 => vga_com_tile_module_n_710, ZN => vga_com_tile_module_n_805);
  vga_com_tile_module_g47930 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_712, A2 => vga_com_tile_module_n_344, B1 => vga_com_tile_module_n_128, B2 => vga_com_tile_module_n_341, ZN => vga_com_tile_module_n_804);
  vga_com_tile_module_g47931 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_610, A2 => vga_com_tile_module_n_586, A3 => vga_com_tile_module_n_114, A4 => vga_com_tile_module_n_110, ZN => vga_com_tile_module_n_829);
  vga_com_tile_module_g47932 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_605, A2 => vga_com_tile_module_n_545, A3 => vga_com_tile_module_n_349, A4 => vga_com_tile_module_n_105, ZN => vga_com_tile_module_n_828);
  vga_com_tile_module_g47933 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_622, A2 => vga_com_tile_module_n_600, A3 => vga_com_tile_module_n_626, A4 => vga_com_tile_module_n_399, ZN => vga_com_tile_module_n_827);
  vga_com_tile_module_g47934 : INVD0BWP7T port map(I => vga_com_tile_module_n_802, ZN => vga_com_tile_module_n_803);
  vga_com_tile_module_g47935 : AOI221D0BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_tile_module_n_569, B1 => vga_com_tile_module_n_425, B2 => vga_com_tile_module_n_50, C => vga_com_tile_module_n_219, ZN => vga_com_tile_module_n_796);
  vga_com_tile_module_g47936 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_48, A2 => vga_com_tile_module_n_572, A3 => vga_com_tile_module_n_425, A4 => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_795);
  vga_com_tile_module_g47937 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_655, A2 => vga_com_tile_module_n_10, B => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_794);
  vga_com_tile_module_g47938 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_169, B1 => vga_com_tile_module_n_712, ZN => vga_com_tile_module_n_793);
  vga_com_tile_module_g47939 : OAI211D1BWP7T port map(A1 => FE_OFN4_vga_com_row_2, A2 => vga_com_tile_module_n_563, B => vga_com_tile_module_n_485, C => vga_com_tile_module_n_302, ZN => vga_com_tile_module_n_792);
  vga_com_tile_module_g47940 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_618, A2 => vga_com_tile_module_n_305, A3 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_791);
  vga_com_tile_module_g47941 : OAI31D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_430, A3 => vga_com_tile_module_n_535, B => vga_com_tile_module_n_495, ZN => vga_com_tile_module_n_790);
  vga_com_tile_module_g47942 : AN3D0BWP7T port map(A1 => vga_com_tile_module_n_630, A2 => vga_com_tile_module_n_506, A3 => vga_com_tile_module_n_114, Z => vga_com_tile_module_n_789);
  vga_com_tile_module_g47943 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_595, A2 => vga_com_tile_module_n_473, B => vga_com_tile_module_n_86, ZN => vga_com_tile_module_n_788);
  vga_com_tile_module_g47944 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_487, A2 => vga_com_tile_module_n_589, A3 => vga_com_tile_module_n_465, ZN => vga_com_tile_module_n_787);
  vga_com_tile_module_g47945 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_661, A2 => vga_com_tile_module_n_583, A3 => vga_com_tile_module_n_301, A4 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_786);
  vga_com_tile_module_g47946 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_123, A2 => vga_com_tile_module_n_178, B => vga_com_tile_module_n_625, C => vga_com_tile_module_n_137, Z => vga_com_tile_module_n_785);
  vga_com_tile_module_g47947 : AOI211D0BWP7T port map(A1 => vga_com_tile_module_n_568, A2 => vga_com_tile_module_n_316, B => vga_com_tile_module_n_199, C => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_784);
  vga_com_tile_module_g47948 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_155, A2 => vga_com_tile_module_n_346, B1 => vga_com_tile_module_n_220, B2 => vga_com_tile_module_n_38, C => vga_com_tile_module_n_681, ZN => vga_com_tile_module_n_783);
  vga_com_tile_module_g47949 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_537, A2 => vga_com_tile_module_n_181, B1 => vga_com_tile_module_n_323, B2 => FE_OFN4_vga_com_row_2, C => vga_com_tile_module_n_106, ZN => vga_com_tile_module_n_782);
  vga_com_tile_module_g47950 : AO221D0BWP7T port map(A1 => vga_com_tile_module_n_22, A2 => vga_com_tile_module_n_570, B1 => vga_com_tile_module_n_25, B2 => vga_com_tile_module_n_11, C => vga_com_tile_module_n_578, Z => vga_com_tile_module_n_781);
  vga_com_tile_module_g47951 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_17, A2 => vga_com_tile_module_n_11, B => vga_com_tile_module_n_596, C => vga_com_tile_module_n_541, ZN => vga_com_tile_module_n_780);
  vga_com_tile_module_g47952 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_632, A2 => vga_com_tile_module_n_544, B1 => vga_com_tile_module_n_378, B2 => vga_com_tile_module_n_110, C1 => vga_com_tile_module_n_377, C2 => vga_com_tile_module_n_105, ZN => vga_com_tile_module_n_779);
  vga_com_tile_module_g47953 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_23, A2 => vga_com_tile_module_n_193, B => vga_com_tile_module_n_696, C => vga_com_tile_module_n_529, ZN => vga_com_tile_module_n_778);
  vga_com_tile_module_g47954 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_585, A2 => vga_com_tile_module_n_448, B1 => vga_com_tile_module_n_16, B2 => vga_com_tile_module_n_321, C => vga_com_tile_module_n_434, ZN => vga_com_tile_module_n_802);
  vga_com_tile_module_g47955 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_714, A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_801);
  vga_com_tile_module_g47956 : AN3D1BWP7T port map(A1 => vga_com_tile_module_n_614, A2 => vga_com_tile_module_n_588, A3 => vga_com_tile_module_n_434, Z => vga_com_tile_module_n_800);
  vga_com_tile_module_g47957 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_591, A2 => vga_com_tile_module_n_371, A3 => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_799);
  vga_com_tile_module_g47958 : ND4D0BWP7T port map(A1 => vga_com_tile_module_n_628, A2 => vga_com_tile_module_n_496, A3 => vga_com_tile_module_n_449, A4 => vga_com_tile_module_n_475, ZN => vga_com_tile_module_n_798);
  vga_com_tile_module_g47959 : CKND2D0BWP7T port map(A1 => vga_com_tile_module_n_748, A2 => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_797);
  vga_com_tile_module_g47960 : INVD0BWP7T port map(I => vga_com_tile_module_n_774, ZN => vga_com_tile_module_n_775);
  vga_com_tile_module_g47961 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_653, A2 => vga_com_tile_module_n_426, B1 => vga_com_tile_module_n_581, B2 => vga_com_tile_module_n_108, ZN => vga_com_tile_module_n_773);
  vga_com_tile_module_g47962 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_599, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_tile_module_n_308, B2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_772);
  vga_com_tile_module_g47963 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_548, A2 => vga_com_tile_module_n_470, A3 => vga_com_tile_module_n_349, B => vga_com_tile_module_n_71, ZN => vga_com_tile_module_n_771);
  vga_com_tile_module_g47964 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_675, A2 => vga_com_tile_module_n_331, B => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_770);
  vga_com_tile_module_g47965 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_106, A2 => vga_com_tile_module_n_291, A3 => vga_com_tile_module_n_501, B => vga_com_tile_module_n_227, ZN => vga_com_tile_module_n_769);
  vga_com_tile_module_g47966 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_658, A2 => vga_com_tile_module_n_467, B => vga_com_tile_module_n_334, ZN => vga_com_tile_module_n_768);
  vga_com_tile_module_g47967 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_522, A2 => vga_com_tile_module_n_489, A3 => vga_com_tile_module_n_438, B => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_767);
  vga_com_tile_module_g47968 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_566, A2 => vga_com_tile_module_n_519, A3 => vga_com_tile_module_n_302, B => vga_com_tile_module_n_159, ZN => vga_com_tile_module_n_766);
  vga_com_tile_module_g47969 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_635, A2 => vga_com_tile_module_n_439, B => vga_com_tile_address(1), ZN => vga_com_tile_module_n_765);
  vga_com_tile_module_g47970 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_638, A2 => vga_com_tile_module_n_21, B1 => vga_com_tile_module_n_203, B2 => vga_com_tile_module_n_144, ZN => vga_com_tile_module_n_764);
  vga_com_tile_module_g47971 : IAO21D0BWP7T port map(A1 => vga_com_tile_module_n_341, A2 => vga_com_tile_module_n_23, B => vga_com_tile_module_n_687, ZN => vga_com_tile_module_n_763);
  vga_com_tile_module_g47972 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_23, A2 => vga_com_tile_module_n_180, A3 => vga_com_tile_module_n_226, B => vga_com_tile_module_n_742, ZN => vga_com_tile_module_n_762);
  vga_com_tile_module_g47973 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_330, A2 => vga_com_tile_module_n_117, B => vga_com_tile_module_n_612, C => vga_com_tile_module_n_106, ZN => vga_com_tile_module_n_761);
  vga_com_tile_module_g47974 : AOI32D1BWP7T port map(A1 => vga_com_tile_module_n_180, A2 => FE_OFN2_vga_com_tile_address_0, A3 => vga_com_tile_module_n_20, B1 => vga_com_tile_module_n_649, B2 => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_760);
  vga_com_tile_module_g47975 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_43, A2 => vga_com_tile_module_n_0, B1 => vga_com_tile_module_n_60, B2 => vga_com_tile_module_n_651, ZN => vga_com_tile_module_n_759);
  vga_com_tile_module_g47976 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_592, A2 => vga_com_tile_module_n_488, B => vga_com_tile_module_n_214, C => vga_com_tile_module_n_3, Z => vga_com_tile_module_n_758);
  vga_com_tile_module_g47977 : OA222D0BWP7T port map(A1 => vga_com_tile_module_n_576, A2 => vga_com_tile_module_n_9, B1 => vga_com_tile_module_n_53, B2 => vga_com_tile_module_n_353, C1 => vga_com_tile_module_n_56, C2 => vga_com_tile_module_n_337, Z => vga_com_tile_module_n_757);
  vga_com_tile_module_g47978 : OAI33D1BWP7T port map(A1 => vga_com_tile_module_n_37, A2 => vga_com_tile_module_n_500, A3 => vga_com_tile_module_n_517, B1 => vga_com_tile_module_n_252, B2 => vga_com_tile_module_n_38, B3 => vga_com_tile_module_n_560, ZN => vga_com_tile_module_n_756);
  vga_com_tile_module_g47979 : OA32D1BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_tile_module_n_183, A3 => vga_com_tile_module_n_571, B1 => vga_com_tile_module_n_340, B2 => vga_com_tile_module_n_425, Z => vga_com_tile_module_n_755);
  vga_com_tile_module_g47980 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_530, A2 => vga_com_tile_module_n_212, B1 => vga_com_tile_module_n_30, B2 => vga_com_tile_module_n_204, C1 => vga_com_tile_module_n_21, C2 => vga_com_tile_module_n_67, ZN => vga_com_tile_module_n_754);
  vga_com_tile_module_g47981 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_138, A2 => vga_com_tile_module_n_347, B1 => vga_com_tile_module_n_32, B2 => vga_com_tile_module_n_512, C1 => vga_com_tile_module_n_177, C2 => vga_com_tile_module_n_129, ZN => vga_com_tile_module_n_753);
  vga_com_tile_module_g47982 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_585, A2 => vga_com_tile_module_n_339, B1 => vga_com_tile_module_n_18, B2 => vga_com_tile_module_n_219, C1 => vga_com_tile_module_n_92, C2 => vga_com_tile_module_n_170, ZN => vga_com_tile_module_n_752);
  vga_com_tile_module_g47983 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_579, A2 => vga_com_tile_module_n_17, B1 => vga_com_tile_module_n_187, B2 => vga_com_tile_module_n_215, C1 => vga_com_tile_module_n_326, C2 => vga_com_tile_module_n_28, ZN => vga_com_tile_module_n_777);
  vga_com_tile_module_g47984 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_47, A2 => vga_com_tile_module_n_25, B => vga_com_tile_module_n_623, C => vga_com_tile_module_n_468, ZN => vga_com_tile_module_n_776);
  vga_com_tile_module_g47985 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_643, A2 => vga_com_tile_module_n_22, B => vga_com_tile_module_n_34, ZN => vga_com_tile_module_n_774);
  vga_com_tile_module_g47986 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_108, A2 => vga_com_tile_module_n_416, B1 => vga_com_tile_module_n_188, B2 => vga_com_tile_module_n_300, C => vga_com_tile_module_n_453, ZN => vga_com_tile_module_n_745);
  vga_com_tile_module_g47987 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_601, A2 => vga_com_tile_module_n_419, ZN => vga_com_tile_module_n_744);
  vga_com_tile_module_g47988 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_658, B1 => vga_com_tile_module_n_168, ZN => vga_com_tile_module_n_743);
  vga_com_tile_module_g47989 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_10, A2 => vga_com_tile_module_n_668, ZN => vga_com_tile_module_n_742);
  vga_com_tile_module_g47990 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_567, A2 => vga_com_tile_module_n_282, A3 => vga_com_tile_module_n_263, B => vga_com_tile_module_n_483, ZN => vga_com_tile_module_n_741);
  vga_com_tile_module_g47991 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_221, A2 => vga_com_tile_module_n_186, B => vga_com_tile_module_n_539, C => vga_com_tile_module_n_458, ZN => vga_com_tile_module_n_740);
  vga_com_tile_module_g47992 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_414, A2 => vga_com_tile_module_n_272, B => vga_com_tile_module_n_502, C => vga_com_tile_module_n_103, ZN => vga_com_tile_module_n_739);
  vga_com_tile_module_g47993 : CKAN2D1BWP7T port map(A1 => vga_com_tile_module_n_607, A2 => vga_com_tile_module_n_677, Z => vga_com_tile_module_n_738);
  vga_com_tile_module_g47994 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_445, A2 => vga_com_tile_module_n_58, A3 => FE_OFN4_vga_com_row_2, B => vga_com_tile_module_n_482, ZN => vga_com_tile_module_n_737);
  vga_com_tile_module_g47995 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_147, A2 => vga_com_tile_module_n_269, B1 => vga_com_column(2), B2 => vga_com_tile_module_n_155, C => vga_com_tile_module_n_606, ZN => vga_com_tile_module_n_736);
  vga_com_tile_module_g47996 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_270, A2 => vga_com_tile_module_n_30, B1 => vga_com_tile_module_n_21, B2 => vga_com_tile_module_n_193, C => vga_com_tile_module_n_659, ZN => vga_com_tile_module_n_735);
  vga_com_tile_module_g47997 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_288, A2 => vga_com_tile_module_n_23, B1 => vga_com_tile_module_n_21, B2 => vga_com_tile_module_n_210, C => vga_com_tile_module_n_661, ZN => vga_com_tile_module_n_734);
  vga_com_tile_module_g47998 : AO221D0BWP7T port map(A1 => vga_com_tile_module_n_472, A2 => vga_com_tile_module_n_10, B1 => vga_com_tile_module_n_25, B2 => vga_com_tile_module_n_81, C => vga_com_tile_module_n_167, Z => vga_com_tile_module_n_733);
  vga_com_tile_module_g47999 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_424, A2 => vga_com_tile_module_n_116, B => vga_com_tile_module_n_62, C => vga_com_tile_module_n_24, ZN => vga_com_tile_module_n_732);
  vga_com_tile_module_g48000 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_412, A2 => vga_com_tile_module_n_38, B1 => vga_com_tile_module_n_63, B2 => vga_com_tile_module_n_37, C => vga_com_tile_module_n_509, ZN => vga_com_tile_module_n_731);
  vga_com_tile_module_g48001 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_322, A2 => vga_com_tile_module_n_25, B1 => vga_com_tile_module_n_243, B2 => vga_com_tile_module_n_20, C => vga_com_tile_module_n_664, ZN => vga_com_tile_module_n_730);
  vga_com_tile_module_g48002 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_447, A2 => vga_com_tile_module_n_16, B1 => vga_com_tile_module_n_12, B2 => vga_com_tile_module_n_61, C => vga_com_tile_module_n_508, ZN => vga_com_tile_module_n_729);
  vga_com_tile_module_g48003 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_120, A2 => vga_com_tile_module_n_186, B1 => vga_com_tile_module_n_16, B2 => vga_com_tile_module_n_340, C => vga_com_tile_module_n_590, ZN => vga_com_tile_module_n_728);
  vga_com_tile_module_g48004 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_571, A2 => vga_com_tile_module_n_447, B => vga_com_tile_module_n_208, ZN => vga_com_tile_module_n_727);
  vga_com_tile_module_g48005 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_303, A2 => vga_com_tile_module_n_278, B1 => vga_com_tile_module_n_441, B2 => vga_com_tile_module_n_34, C => vga_com_tile_module_n_598, ZN => vga_com_tile_module_n_726);
  vga_com_tile_module_g48006 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_431, A2 => vga_com_tile_module_n_18, B1 => vga_com_tile_module_n_16, B2 => vga_com_tile_module_n_357, C => vga_com_tile_module_n_511, ZN => vga_com_tile_module_n_725);
  vga_com_tile_module_g48007 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_436, A2 => vga_com_tile_module_n_427, B1 => vga_com_tile_module_n_16, B2 => vga_com_tile_module_n_261, C => vga_com_tile_module_n_514, ZN => vga_com_tile_module_n_724);
  vga_com_tile_module_g48008 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_401, A2 => vga_com_tile_module_n_222, B1 => vga_com_tile_module_n_78, B2 => vga_com_tile_module_n_112, C => vga_com_tile_module_n_497, ZN => vga_com_tile_module_n_723);
  vga_com_tile_module_g48009 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_455, A2 => vga_com_tile_module_n_16, B1 => vga_com_tile_module_n_104, B2 => vga_com_tile_module_n_191, C => vga_com_tile_module_n_376, ZN => vga_com_tile_module_n_722);
  vga_com_tile_module_g48010 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_416, A2 => vga_com_tile_module_n_203, B1 => vga_com_tile_module_n_142, B2 => vga_com_tile_module_n_350, C => vga_com_tile_module_n_494, ZN => vga_com_tile_module_n_721);
  vga_com_tile_module_g48011 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_356, A2 => vga_com_tile_module_n_30, B => vga_com_tile_module_n_671, ZN => vga_com_tile_module_n_720);
  vga_com_tile_module_g48012 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_552, A2 => vga_com_column(2), B => vga_com_tile_module_n_436, ZN => vga_com_tile_module_n_719);
  vga_com_tile_module_g48013 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_567, A2 => vga_com_tile_module_n_12, B => vga_com_tile_module_n_238, ZN => vga_com_tile_module_n_718);
  vga_com_tile_module_g48014 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_18, A2 => vga_com_tile_module_n_415, B => vga_com_tile_module_n_617, C => vga_com_tile_module_n_449, ZN => vga_com_tile_module_n_717);
  vga_com_tile_module_g48015 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_16, A2 => vga_com_tile_module_n_11, B1 => vga_com_tile_module_n_114, B2 => vga_com_tile_module_n_223, C => vga_com_tile_module_n_510, ZN => vga_com_tile_module_n_716);
  vga_com_tile_module_g48016 : OAI31D0BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_tile_module_n_317, A3 => vga_com_tile_module_n_427, B => vga_com_tile_module_n_101, ZN => vga_com_tile_module_n_751);
  vga_com_tile_module_g48017 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_362, A2 => vga_com_tile_module_n_171, B => vga_com_tile_module_n_568, C => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_750);
  vga_com_tile_module_g48018 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_667, A2 => vga_com_tile_module_n_22, ZN => vga_com_tile_module_n_749);
  vga_com_tile_module_g48019 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_440, A2 => vga_com_tile_module_n_16, B1 => vga_com_tile_module_n_112, B2 => vga_com_tile_module_n_262, C => vga_com_tile_module_n_575, ZN => vga_com_tile_module_n_748);
  vga_com_tile_module_g48020 : NR4D0BWP7T port map(A1 => vga_com_tile_module_n_490, A2 => vga_com_tile_module_n_398, A3 => vga_com_tile_module_n_293, A4 => vga_com_tile_module_n_465, ZN => vga_com_tile_module_n_747);
  vga_com_tile_module_g48021 : INR2XD0BWP7T port map(A1 => vga_com_tile_module_n_666, B1 => vga_com_tile_module_n_460, ZN => vga_com_tile_module_n_746);
  vga_com_tile_module_g48022 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_526, A2 => vga_com_tile_module_n_26, B1 => vga_com_tile_module_n_357, B2 => vga_com_tile_module_n_29, ZN => vga_com_tile_module_n_711);
  vga_com_tile_module_g48023 : AOI21D0BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_tile_module_n_570, B => vga_com_tile_module_n_178, ZN => vga_com_tile_module_n_710);
  vga_com_tile_module_g48024 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_425, A2 => vga_com_tile_module_n_180, B => vga_com_tile_module_n_269, C => vga_com_tile_module_n_132, ZN => vga_com_tile_module_n_709);
  vga_com_tile_module_g48025 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_139, A2 => vga_com_tile_module_n_11, B => vga_com_tile_module_n_631, ZN => vga_com_tile_module_n_708);
  vga_com_tile_module_g48026 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_203, A2 => vga_com_tile_module_n_216, B => vga_com_tile_module_n_603, C => vga_com_tile_module_n_549, ZN => vga_com_tile_module_n_707);
  vga_com_tile_module_g48027 : OA22D0BWP7T port map(A1 => vga_com_tile_module_n_579, A2 => vga_com_tile_module_n_16, B1 => vga_com_tile_module_n_112, B2 => vga_com_tile_module_n_290, Z => vga_com_tile_module_n_706);
  vga_com_tile_module_g48028 : AN3D1BWP7T port map(A1 => vga_com_tile_module_n_82, A2 => vga_com_tile_module_n_580, A3 => vga_com_tile_module_n_2, Z => vga_com_tile_module_n_705);
  vga_com_tile_module_g48029 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_568, A2 => vga_com_tile_module_n_11, B => vga_com_tile_module_n_76, ZN => vga_com_tile_module_n_704);
  vga_com_tile_module_g48030 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_317, A2 => vga_com_tile_module_n_425, B => vga_com_tile_module_n_198, C => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_703);
  vga_com_tile_module_g48031 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_1060, A2 => vga_com_tile_module_n_9, B1 => vga_com_tile_module_n_562, B2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_702);
  vga_com_tile_module_g48032 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_558, A2 => vga_com_tile_module_n_438, B => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_701);
  vga_com_tile_module_g48033 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_141, A2 => vga_com_tile_module_n_388, B => vga_com_tile_module_n_516, C => vga_com_tile_module_n_195, ZN => vga_com_tile_module_n_700);
  vga_com_tile_module_g48034 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_108, A2 => vga_com_tile_module_n_315, A3 => vga_com_tile_module_n_8, B => vga_com_tile_module_n_621, ZN => vga_com_tile_module_n_699);
  vga_com_tile_module_g48035 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_268, A2 => vga_com_tile_module_n_436, B => vga_com_tile_module_n_652, ZN => vga_com_tile_module_n_698);
  vga_com_tile_module_g48036 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_561, A2 => vga_com_tile_module_n_464, B1 => vga_com_tile_module_n_26, B2 => vga_com_tile_module_n_429, C1 => vga_com_tile_module_n_184, C2 => vga_com_tile_module_n_324, ZN => vga_com_tile_module_n_697);
  vga_com_tile_module_g48037 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_426, A2 => vga_com_tile_module_n_255, B1 => vga_com_tile_module_n_195, B2 => vga_com_tile_module_n_20, C1 => vga_com_tile_module_n_360, C2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_696);
  vga_com_tile_module_g48038 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_1060, A2 => vga_com_tile_module_n_34, B1 => vga_com_tile_module_n_457, B2 => vga_com_tile_module_n_33, ZN => vga_com_tile_module_n_695);
  vga_com_tile_module_g48039 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_25, A2 => vga_com_column(0), B => vga_com_tile_module_n_604, ZN => vga_com_tile_module_n_694);
  vga_com_tile_module_g48040 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_382, A2 => vga_com_tile_module_n_275, B1 => vga_com_tile_module_n_63, B2 => vga_com_tile_module_n_21, C1 => vga_com_tile_module_n_30, C2 => vga_com_tile_module_n_224, ZN => vga_com_tile_module_n_693);
  vga_com_tile_module_g48041 : IAO21D0BWP7T port map(A1 => vga_com_tile_module_n_156, A2 => vga_com_tile_module_n_29, B => vga_com_tile_module_n_602, ZN => vga_com_tile_module_n_692);
  vga_com_tile_module_g48042 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_576, A2 => vga_com_tile_module_n_37, B1 => vga_com_tile_module_n_421, B2 => vga_com_tile_module_n_41, ZN => vga_com_tile_module_n_691);
  vga_com_tile_module_g48043 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_20, A2 => vga_com_tile_module_n_574, B1 => vga_com_tile_module_n_181, B2 => vga_com_tile_module_n_31, C1 => vga_com_tile_module_n_209, C2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_690);
  vga_com_tile_module_g48044 : OAI32D1BWP7T port map(A1 => vga_com_tile_module_n_46, A2 => vga_com_tile_module_n_266, A3 => vga_com_tile_module_n_427, B1 => vga_com_tile_module_n_50, B2 => vga_com_tile_module_n_73, ZN => vga_com_tile_module_n_689);
  vga_com_tile_module_g48045 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_308, A2 => vga_com_tile_module_n_32, B1 => vga_com_tile_module_n_432, B2 => vga_com_tile_module_n_107, C1 => vga_com_tile_module_n_310, C2 => vga_com_tile_module_n_189, ZN => vga_com_tile_module_n_688);
  vga_com_tile_module_g48046 : AOI32D0BWP7T port map(A1 => vga_com_tile_module_n_450, A2 => vga_com_tile_module_n_277, A3 => vga_com_tile_module_n_188, B1 => vga_com_tile_module_n_108, B2 => vga_com_tile_module_n_121, ZN => vga_com_tile_module_n_687);
  vga_com_tile_module_g48047 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_577, A2 => vga_com_tile_module_n_107, B1 => vga_com_tile_module_n_584, B2 => vga_com_tile_module_n_189, ZN => vga_com_tile_module_n_686);
  vga_com_tile_module_g48048 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_112, A2 => vga_com_tile_module_n_88, B1 => vga_com_tile_module_n_555, B2 => vga_com_tile_module_n_73, ZN => vga_com_tile_module_n_685);
  vga_com_tile_module_g48049 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_276, A2 => vga_com_tile_module_n_28, B => vga_com_tile_module_n_532, C => vga_com_tile_module_n_379, ZN => vga_com_tile_module_n_684);
  vga_com_tile_module_g48050 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_528, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_151, B2 => vga_com_tile_module_n_455, ZN => vga_com_tile_module_n_683);
  vga_com_tile_module_g48051 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_581, A2 => vga_com_tile_module_n_19, B1 => vga_com_tile_module_n_300, B2 => vga_com_tile_module_n_29, ZN => vga_com_tile_module_n_682);
  vga_com_tile_module_g48052 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_525, A2 => vga_com_tile_module_n_188, B1 => vga_com_tile_module_n_149, B2 => vga_com_tile_module_n_232, ZN => vga_com_tile_module_n_681);
  vga_com_tile_module_g48053 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_476, A2 => vga_com_tile_module_n_2, B1 => vga_com_tile_module_n_543, B2 => vga_com_tile_module_n_37, ZN => vga_com_tile_module_n_680);
  vga_com_tile_module_g48054 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_546, A2 => vga_com_tile_module_n_209, B1 => vga_com_tile_module_n_106, B2 => vga_com_tile_module_n_210, ZN => vga_com_tile_module_n_679);
  vga_com_tile_module_g48055 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_412, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_tile_module_n_9, B2 => vga_com_tile_module_n_63, C1 => vga_com_tile_module_n_58, C2 => vga_com_tile_module_n_29, ZN => vga_com_tile_module_n_715);
  vga_com_tile_module_g48056 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_551, A2 => vga_com_tile_module_n_261, B1 => vga_com_tile_module_n_326, B2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_714);
  vga_com_tile_module_g48057 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_326, A2 => FE_OFN3_vga_com_row_1, B => vga_com_tile_module_n_582, C => vga_com_tile_module_n_37, Z => vga_com_tile_module_n_713);
  vga_com_tile_module_g48058 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_568, A2 => vga_com_tile_module_n_178, B => vga_com_tile_module_n_62, ZN => vga_com_tile_module_n_712);
  vga_com_tile_module_g48059 : CKND1BWP7T port map(I => vga_com_tile_module_n_673, ZN => vga_com_tile_module_n_674);
  vga_com_tile_module_g48060 : INVD0BWP7T port map(I => vga_com_tile_module_n_659, ZN => vga_com_tile_module_n_660);
  vga_com_tile_module_g48061 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_568, A2 => vga_com_tile_module_n_570, ZN => vga_com_tile_module_n_657);
  vga_com_tile_module_g48062 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_404, A2 => vga_com_tile_module_n_58, B => vga_com_tile_module_n_390, Z => vga_com_tile_module_n_656);
  vga_com_tile_module_g48063 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_567, A2 => vga_com_tile_module_n_65, ZN => vga_com_tile_module_n_655);
  vga_com_tile_module_g48064 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_572, A2 => vga_com_tile_module_n_427, ZN => vga_com_tile_module_n_654);
  vga_com_tile_module_g48065 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_102, A2 => vga_com_tile_module_n_35, B => vga_com_tile_module_n_380, C => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_653);
  vga_com_tile_module_g48066 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_146, A2 => vga_com_tile_module_n_235, B1 => vga_com_tile_module_n_16, B2 => vga_com_tile_module_n_260, C => vga_com_tile_module_n_434, ZN => vga_com_tile_module_n_652);
  vga_com_tile_module_g48067 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_332, A2 => vga_com_tile_module_n_22, B1 => vga_com_tile_module_n_324, B2 => vga_com_tile_module_n_25, C => vga_com_tile_module_n_414, ZN => vga_com_tile_module_n_651);
  vga_com_tile_module_g48068 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_359, A2 => FE_OFN3_vga_com_row_1, B1 => vga_com_tile_module_n_182, B2 => vga_com_tile_module_n_20, C => vga_com_tile_module_n_167, ZN => vga_com_tile_module_n_650);
  vga_com_tile_module_g48069 : AO221D0BWP7T port map(A1 => vga_com_tile_module_n_294, A2 => vga_com_tile_module_n_66, B1 => vga_com_tile_module_n_191, B2 => vga_com_tile_module_n_103, C => vga_com_tile_module_n_352, Z => vga_com_tile_module_n_649);
  vga_com_tile_module_g48070 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_276, A2 => FE_OFN3_vga_com_row_1, B1 => vga_com_tile_module_n_53, B2 => vga_com_tile_module_n_226, C => vga_com_tile_module_n_405, ZN => vga_com_tile_module_n_648);
  vga_com_tile_module_g48071 : OA221D0BWP7T port map(A1 => vga_com_tile_module_n_342, A2 => FE_OFN4_vga_com_row_2, B1 => vga_com_tile_module_n_10, B2 => vga_com_tile_module_n_333, C => vga_com_tile_module_n_184, Z => vga_com_tile_module_n_647);
  vga_com_tile_module_g48072 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_355, A2 => vga_com_tile_module_n_106, B1 => vga_com_tile_module_n_109, B2 => vga_com_tile_module_n_79, C => vga_com_tile_module_n_504, ZN => vga_com_tile_module_n_646);
  vga_com_tile_module_g48073 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_183, A2 => vga_com_tile_module_n_137, B1 => vga_com_tile_module_n_188, B2 => vga_com_tile_module_n_192, C => vga_com_tile_module_n_491, ZN => vga_com_tile_module_n_645);
  vga_com_tile_module_g48074 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_355, A2 => vga_com_tile_module_n_22, B1 => vga_com_tile_module_n_163, B2 => vga_com_tile_module_n_20, C => vga_com_tile_module_n_493, ZN => vga_com_tile_module_n_644);
  vga_com_tile_module_g48075 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_446, A2 => FE_OFN3_vga_com_row_1, B => vga_com_tile_module_n_582, ZN => vga_com_tile_module_n_643);
  vga_com_tile_module_g48076 : OAI31D0BWP7T port map(A1 => vga_com_tile_module_n_178, A2 => vga_com_tile_module_n_106, A3 => vga_com_tile_module_n_257, B => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_642);
  vga_com_tile_module_g48077 : AOI31D0BWP7T port map(A1 => vga_com_tile_module_n_120, A2 => vga_com_tile_module_n_47, A3 => vga_com_tile_module_n_20, B => vga_com_tile_module_n_503, ZN => vga_com_tile_module_n_641);
  vga_com_tile_module_g48078 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_18, A2 => vga_com_tile_module_n_261, B => vga_com_tile_module_n_403, C => vga_com_tile_module_n_407, ZN => vga_com_tile_module_n_640);
  vga_com_tile_module_g48079 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_145, A2 => vga_com_tile_module_n_181, B => vga_com_tile_module_n_575, ZN => vga_com_tile_module_n_639);
  vga_com_tile_module_g48080 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_471, A2 => vga_com_tile_module_n_38, A3 => vga_com_tile_module_n_173, ZN => vga_com_tile_module_n_638);
  vga_com_tile_module_g48081 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_323, A2 => vga_com_tile_module_n_348, B => vga_com_tile_module_n_433, C => vga_com_tile_module_n_291, ZN => vga_com_tile_module_n_637);
  vga_com_tile_module_g48082 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_422, A2 => vga_com_tile_module_n_18, B1 => vga_com_tile_module_n_329, B2 => vga_com_tile_module_n_29, ZN => vga_com_tile_module_n_636);
  vga_com_tile_module_g48083 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_29, A2 => vga_com_tile_module_n_259, B => vga_com_tile_module_n_463, C => vga_com_tile_module_n_299, ZN => vga_com_tile_module_n_635);
  vga_com_tile_module_g48084 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_168, A2 => vga_com_tile_module_n_25, B => vga_com_tile_module_n_400, C => vga_com_tile_module_n_461, ZN => vga_com_tile_module_n_634);
  vga_com_tile_module_g48085 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_424, A2 => vga_com_tile_module_n_246, B => vga_com_tile_module_n_175, ZN => vga_com_tile_module_n_633);
  vga_com_tile_module_g48086 : AN3D0BWP7T port map(A1 => vga_com_tile_module_n_450, A2 => vga_com_tile_module_n_179, A3 => FE_OFN3_vga_com_row_1, Z => vga_com_tile_module_n_632);
  vga_com_tile_module_g48087 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_282, A2 => vga_com_tile_module_n_265, B => vga_com_tile_module_n_381, C => vga_com_tile_module_n_477, Z => vga_com_tile_module_n_631);
  vga_com_tile_module_g48088 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_573, B1 => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_678);
  vga_com_tile_module_g48089 : AO221D0BWP7T port map(A1 => vga_com_tile_module_n_341, A2 => FE_OFN1_vga_com_row_0, B1 => vga_com_tile_module_n_164, B2 => vga_com_tile_module_n_8, C => vga_com_tile_module_n_18, Z => vga_com_tile_module_n_677);
  vga_com_tile_module_g48090 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_332, A2 => FE_OFN1_vga_com_row_0, B1 => vga_com_tile_module_n_8, B2 => vga_com_tile_module_n_88, C => vga_com_tile_module_n_364, ZN => vga_com_tile_module_n_676);
  vga_com_tile_module_g48091 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_568, A2 => vga_com_tile_module_n_195, ZN => vga_com_tile_module_n_675);
  vga_com_tile_module_g48092 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_435, A2 => vga_com_tile_module_n_20, B => vga_com_tile_module_n_298, ZN => vga_com_tile_module_n_673);
  vga_com_tile_module_g48093 : AOI221D1BWP7T port map(A1 => vga_com_tile_module_n_280, A2 => vga_com_tile_module_n_25, B1 => vga_com_tile_module_n_221, B2 => vga_com_tile_module_n_22, C => vga_com_tile_module_n_309, ZN => vga_com_tile_module_n_672);
  vga_com_tile_module_g48094 : AOI221D1BWP7T port map(A1 => vga_com_tile_module_n_314, A2 => FE_OFN3_vga_com_row_1, B1 => vga_com_tile_module_n_120, B2 => vga_com_tile_module_n_20, C => vga_com_tile_module_n_22, ZN => vga_com_tile_module_n_671);
  vga_com_tile_module_g48095 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_265, A2 => vga_com_tile_module_n_22, B1 => vga_com_tile_module_n_193, B2 => vga_com_tile_module_n_25, C => vga_com_tile_module_n_178, ZN => vga_com_tile_module_n_670);
  vga_com_tile_module_g48096 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_567, A2 => vga_com_tile_module_n_192, ZN => vga_com_tile_module_n_669);
  vga_com_tile_module_g48097 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_261, A2 => vga_com_tile_module_n_574, ZN => vga_com_tile_module_n_668);
  vga_com_tile_module_g48098 : CKAN2D1BWP7T port map(A1 => vga_com_tile_module_n_584, A2 => vga_com_tile_module_n_11, Z => vga_com_tile_module_n_667);
  vga_com_tile_module_g48099 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_387, A2 => FE_OFN3_vga_com_row_1, B => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_666);
  vga_com_tile_module_g48100 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_572, B1 => vga_com_tile_module_n_43, ZN => vga_com_tile_module_n_665);
  vga_com_tile_module_g48101 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_315, A2 => vga_com_tile_module_n_30, B => vga_com_tile_module_n_583, ZN => vga_com_tile_module_n_664);
  vga_com_tile_module_g48102 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_553, A2 => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_663);
  vga_com_tile_module_g48103 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_420, A2 => vga_com_tile_module_n_16, B1 => vga_com_tile_module_n_277, B2 => vga_com_tile_module_n_26, ZN => vga_com_tile_module_n_662);
  vga_com_tile_module_g48104 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_428, A2 => vga_com_tile_module_n_31, B1 => vga_com_tile_module_n_225, B2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_661);
  vga_com_tile_module_g48105 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_567, A2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_659);
  vga_com_tile_module_g48106 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_568, A2 => vga_com_tile_module_n_179, ZN => vga_com_tile_module_n_658);
  vga_com_tile_module_g48107 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_451, A2 => vga_com_tile_module_n_28, B1 => vga_com_tile_module_n_320, B2 => vga_com_tile_module_n_117, C1 => vga_com_tile_module_n_181, C2 => vga_com_tile_module_n_103, ZN => vga_com_tile_module_n_628);
  vga_com_tile_module_g48108 : OAI211D0BWP7T port map(A1 => vga_com_tile_module_n_8, A2 => vga_com_tile_module_n_345, B => vga_com_tile_module_n_298, C => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_627);
  vga_com_tile_module_g48109 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_430, A2 => vga_com_tile_module_n_319, B => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_626);
  vga_com_tile_module_g48110 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_411, A2 => vga_com_tile_module_n_321, B1 => vga_com_tile_module_n_189, B2 => vga_com_tile_module_n_272, ZN => vga_com_tile_module_n_625);
  vga_com_tile_module_g48111 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_53, A2 => vga_com_tile_module_n_201, B => vga_com_tile_module_n_481, C => vga_com_tile_module_n_459, ZN => vga_com_tile_module_n_624);
  vga_com_tile_module_g48112 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_462, A2 => vga_com_tile_module_n_30, B => vga_com_tile_module_n_209, ZN => vga_com_tile_module_n_623);
  vga_com_tile_module_g48113 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_428, A2 => vga_com_tile_module_n_113, B1 => vga_com_tile_module_n_454, B2 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_622);
  vga_com_tile_module_g48114 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_445, A2 => vga_com_tile_module_n_189, B1 => vga_com_tile_module_n_250, B2 => vga_com_tile_module_n_73, ZN => vga_com_tile_module_n_621);
  vga_com_tile_module_g48115 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_166, A2 => vga_com_tile_module_n_245, B => vga_com_tile_module_n_253, C => vga_com_tile_module_n_394, ZN => vga_com_tile_module_n_620);
  vga_com_tile_module_g48116 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_277, A2 => vga_com_tile_module_n_152, B => vga_com_tile_module_n_396, C => vga_com_tile_module_n_372, ZN => vga_com_tile_module_n_619);
  vga_com_tile_module_g48117 : OAI211D1BWP7T port map(A1 => vga_com_tile_module_n_199, A2 => vga_com_tile_module_n_184, B => vga_com_tile_module_n_373, C => vga_com_tile_module_n_375, ZN => vga_com_tile_module_n_618);
  vga_com_tile_module_g48118 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_371, A2 => vga_com_tile_module_n_29, B => vga_com_tile_module_n_540, Z => vga_com_tile_module_n_617);
  vga_com_tile_module_g48119 : OA222D0BWP7T port map(A1 => vga_com_tile_module_n_424, A2 => vga_com_tile_module_n_436, B1 => vga_com_tile_module_n_118, B2 => vga_com_tile_module_n_120, C1 => vga_com_tile_module_n_190, C2 => vga_com_tile_module_n_146, Z => vga_com_tile_module_n_616);
  vga_com_tile_module_g48120 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_469, A2 => vga_com_tile_module_n_8, B => vga_com_tile_module_n_515, ZN => vga_com_tile_module_n_615);
  vga_com_tile_module_g48121 : OA222D0BWP7T port map(A1 => vga_com_tile_module_n_444, A2 => vga_com_tile_module_n_339, B1 => vga_com_tile_module_n_118, B2 => vga_com_tile_module_n_360, C1 => vga_com_tile_module_n_104, C2 => vga_com_tile_module_n_328, Z => vga_com_tile_module_n_614);
  vga_com_tile_module_g48122 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_134, A2 => vga_com_tile_module_n_244, B => vga_com_tile_module_n_505, ZN => vga_com_tile_module_n_613);
  vga_com_tile_module_g48123 : AO222D0BWP7T port map(A1 => vga_com_tile_module_n_341, A2 => vga_com_tile_module_n_19, B1 => vga_com_tile_module_n_393, B2 => vga_com_tile_module_n_58, C1 => vga_com_tile_module_n_365, C2 => vga_com_tile_module_n_27, Z => vga_com_tile_module_n_612);
  vga_com_tile_module_g48124 : OA221D0BWP7T port map(A1 => vga_com_tile_module_n_194, A2 => vga_com_tile_module_n_23, B1 => vga_com_tile_module_n_24, B2 => vga_com_tile_module_n_226, C => vga_com_tile_module_n_389, Z => vga_com_tile_module_n_611);
  vga_com_tile_module_g48125 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_446, A2 => vga_com_tile_module_n_57, B => vga_com_tile_module_n_498, ZN => vga_com_tile_module_n_610);
  vga_com_tile_module_g48126 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_206, A2 => vga_com_tile_module_n_25, B1 => vga_com_tile_module_n_454, B2 => vga_com_tile_module_n_10, C => vga_com_tile_module_n_468, ZN => vga_com_tile_module_n_609);
  vga_com_tile_module_g48127 : OAI222D0BWP7T port map(A1 => vga_com_tile_module_n_149, A2 => vga_com_tile_module_n_330, B1 => vga_com_tile_module_n_213, B2 => vga_com_tile_module_n_165, C1 => vga_com_tile_module_n_73, C2 => vga_com_tile_module_n_134, ZN => vga_com_tile_module_n_608);
  vga_com_tile_module_g48128 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_356, A2 => vga_com_tile_module_n_103, B1 => vga_com_tile_module_n_322, B2 => vga_com_tile_module_n_185, C1 => vga_com_tile_module_n_187, C2 => vga_com_tile_module_n_244, ZN => vga_com_tile_module_n_607);
  vga_com_tile_module_g48129 : AOI32D1BWP7T port map(A1 => vga_com_tile_module_n_279, A2 => vga_com_tile_module_n_39, A3 => vga_com_tile_module_n_20, B1 => vga_com_tile_module_n_133, B2 => vga_com_tile_module_n_194, ZN => vga_com_tile_module_n_606);
  vga_com_tile_module_g48130 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_423, A2 => vga_com_tile_module_n_316, B1 => vga_com_tile_module_n_185, B2 => vga_com_tile_module_n_161, ZN => vga_com_tile_module_n_605);
  vga_com_tile_module_g48131 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_418, A2 => FE_OFN3_vga_com_row_1, B1 => vga_com_tile_module_n_23, B2 => vga_com_tile_module_n_75, ZN => vga_com_tile_module_n_604);
  vga_com_tile_module_g48132 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_446, A2 => vga_com_tile_module_n_354, B1 => vga_com_tile_module_n_136, B2 => vga_com_tile_module_n_179, ZN => vga_com_tile_module_n_603);
  vga_com_tile_module_g48133 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_197, A2 => vga_com_tile_module_n_104, B1 => vga_com_tile_module_n_409, B2 => vga_com_tile_module_n_443, ZN => vga_com_tile_module_n_602);
  vga_com_tile_module_g48134 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_221, A2 => vga_com_tile_module_n_20, B => vga_com_tile_module_n_383, C => vga_com_tile_module_n_254, ZN => vga_com_tile_module_n_601);
  vga_com_tile_module_g48135 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_437, A2 => vga_com_tile_module_n_27, B1 => vga_com_tile_module_n_186, B2 => vga_com_tile_module_n_324, ZN => vga_com_tile_module_n_600);
  vga_com_tile_module_g48136 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_431, A2 => vga_com_tile_module_n_10, B1 => vga_com_tile_module_n_287, B2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_599);
  vga_com_tile_module_g48137 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_469, A2 => vga_com_tile_module_n_20, B1 => vga_com_tile_module_n_125, B2 => vga_com_tile_module_n_262, ZN => vga_com_tile_module_n_598);
  vga_com_tile_module_g48138 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_441, A2 => vga_com_tile_module_n_123, B1 => vga_com_tile_module_n_344, B2 => vga_com_tile_module_n_316, ZN => vga_com_tile_module_n_597);
  vga_com_tile_module_g48139 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_437, A2 => vga_com_tile_module_n_18, B1 => vga_com_tile_module_n_294, B2 => vga_com_tile_module_n_85, ZN => vga_com_tile_module_n_596);
  vga_com_tile_module_g48140 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_107, A2 => vga_com_tile_module_n_415, B1 => vga_com_tile_module_n_188, B2 => vga_com_tile_module_n_342, ZN => vga_com_tile_module_n_595);
  vga_com_tile_module_g48141 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_447, A2 => vga_com_tile_module_n_27, B1 => vga_com_tile_module_n_187, B2 => vga_com_tile_module_n_200, ZN => vga_com_tile_module_n_594);
  vga_com_tile_module_g48142 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_448, A2 => vga_com_tile_module_n_134, B1 => vga_com_tile_module_n_141, B2 => vga_com_tile_module_n_199, ZN => vga_com_tile_module_n_593);
  vga_com_tile_module_g48143 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_321, A2 => vga_com_tile_module_n_142, B1 => vga_com_tile_module_n_412, B2 => vga_com_tile_module_n_126, ZN => vga_com_tile_module_n_592);
  vga_com_tile_module_g48144 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_315, A2 => vga_com_tile_module_n_61, B1 => vga_com_tile_module_n_445, B2 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_591);
  vga_com_tile_module_g48145 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_467, A2 => vga_com_tile_module_n_103, B1 => vga_com_tile_module_n_329, B2 => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_590);
  vga_com_tile_module_g48146 : AO22D0BWP7T port map(A1 => vga_com_tile_module_n_428, A2 => vga_com_tile_module_n_28, B1 => vga_com_tile_module_n_78, B2 => vga_com_tile_module_n_174, Z => vga_com_tile_module_n_589);
  vga_com_tile_module_g48147 : OA22D0BWP7T port map(A1 => vga_com_tile_module_n_428, A2 => vga_com_tile_module_n_110, B1 => vga_com_tile_module_n_186, B2 => vga_com_tile_module_n_290, Z => vga_com_tile_module_n_588);
  vga_com_tile_module_g48148 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_452, A2 => vga_com_tile_module_n_135, B1 => vga_com_tile_module_n_366, B2 => vga_com_tile_module_n_334, ZN => vga_com_tile_module_n_587);
  vga_com_tile_module_g48149 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_428, A2 => vga_com_tile_module_n_187, B1 => vga_com_tile_module_n_27, B2 => vga_com_tile_module_n_78, ZN => vga_com_tile_module_n_586);
  vga_com_tile_module_g48150 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_392, A2 => vga_com_tile_module_n_121, B1 => vga_com_tile_module_n_314, B2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_630);
  vga_com_tile_module_g48151 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_408, A2 => vga_com_tile_module_n_29, B1 => vga_com_tile_module_n_286, B2 => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_629);
  vga_com_tile_module_g48153 : INVD0BWP7T port map(I => vga_com_tile_module_n_569, ZN => vga_com_tile_module_n_570);
  vga_com_tile_module_g48154 : INVD1BWP7T port map(I => vga_com_tile_module_n_568, ZN => vga_com_tile_module_n_567);
  vga_com_tile_module_g48155 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_258, A2 => vga_com_tile_module_n_57, B1 => vga_com_tile_module_n_199, B2 => vga_com_tile_module_n_52, C1 => vga_com_tile_module_n_19, C2 => vga_com_tile_module_n_207, ZN => vga_com_tile_module_n_566);
  vga_com_tile_module_g48156 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_427, A2 => vga_com_tile_module_n_119, ZN => vga_com_tile_module_n_565);
  vga_com_tile_module_g48157 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_466, B1 => vga_com_tile_module_n_203, ZN => vga_com_tile_module_n_564);
  vga_com_tile_module_g48158 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_333, B1 => vga_com_tile_module_n_429, ZN => vga_com_tile_module_n_563);
  vga_com_tile_module_g48159 : CKAN2D1BWP7T port map(A1 => vga_com_tile_module_n_457, A2 => vga_com_tile_module_n_121, Z => vga_com_tile_module_n_562);
  vga_com_tile_module_g48160 : OAI32D1BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_tile_module_n_204, A3 => vga_com_tile_module_n_183, B1 => FE_OFN3_vga_com_row_1, B2 => vga_com_tile_module_n_327, ZN => vga_com_tile_module_n_561);
  vga_com_tile_module_g48161 : OAI32D1BWP7T port map(A1 => vga_com_tile_module_n_24, A2 => vga_com_tile_module_n_74, A3 => vga_com_tile_module_n_200, B1 => vga_com_tile_module_n_21, B2 => vga_com_tile_module_n_265, ZN => vga_com_tile_module_n_560);
  vga_com_tile_module_g48162 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_413, B1 => vga_com_tile_module_n_397, ZN => vga_com_tile_module_n_559);
  vga_com_tile_module_g48163 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_197, A2 => vga_com_tile_module_n_113, B1 => vga_com_tile_module_n_185, B2 => vga_com_tile_module_n_80, C => vga_com_tile_module_n_460, ZN => vga_com_tile_module_n_558);
  vga_com_tile_module_g48164 : AOI221D0BWP7T port map(A1 => vga_com_tile_module_n_109, A2 => vga_com_column(1), B1 => FE_OFN4_vga_com_row_2, B2 => vga_com_tile_module_n_4, C => vga_com_tile_module_n_374, ZN => vga_com_tile_module_n_557);
  vga_com_tile_module_g48165 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_311, A2 => vga_com_tile_module_n_147, B1 => vga_com_tile_module_n_153, B2 => vga_com_tile_module_n_238, ZN => vga_com_tile_module_n_556);
  vga_com_tile_module_g48166 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_266, A2 => vga_com_column(1), B => vga_com_tile_module_n_458, ZN => vga_com_tile_module_n_555);
  vga_com_tile_module_g48167 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_273, A2 => FE_OFN3_vga_com_row_1, B => vga_com_tile_module_n_424, ZN => vga_com_tile_module_n_554);
  vga_com_tile_module_g48168 : OAI211D1BWP7T port map(A1 => FE_OFN4_vga_com_row_2, A2 => vga_com_tile_module_n_62, B => vga_com_tile_module_n_307, C => vga_com_tile_module_n_349, ZN => vga_com_tile_module_n_553);
  vga_com_tile_module_g48169 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_309, A2 => vga_com_tile_module_n_296, B => vga_com_tile_module_n_249, Z => vga_com_tile_module_n_552);
  vga_com_tile_module_g48170 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_321, A2 => FE_OFN3_vga_com_row_1, B => vga_com_tile_module_n_30, ZN => vga_com_tile_module_n_551);
  vga_com_tile_module_g48171 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_200, A2 => vga_com_tile_module_n_29, B => vga_com_tile_module_n_463, Z => vga_com_tile_module_n_550);
  vga_com_tile_module_g48172 : IAO21D0BWP7T port map(A1 => vga_com_tile_module_n_34, A2 => vga_com_tile_module_n_348, B => vga_com_tile_module_n_435, ZN => vga_com_tile_module_n_549);
  vga_com_tile_module_g48173 : IND3D1BWP7T port map(A1 => vga_com_tile_module_n_357, B1 => vga_com_tile_module_n_9, B2 => vga_com_tile_module_n_297, ZN => vga_com_tile_module_n_548);
  vga_com_tile_module_g48174 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_361, A2 => vga_com_tile_module_n_31, B1 => vga_com_tile_module_n_167, B2 => vga_com_tile_module_n_75, ZN => vga_com_tile_module_n_547);
  vga_com_tile_module_g48175 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_328, A2 => vga_com_tile_module_n_16, B => vga_com_tile_module_n_118, Z => vga_com_tile_module_n_546);
  vga_com_tile_module_g48176 : OAI211D1BWP7T port map(A1 => FE_OFN3_vga_com_row_1, A2 => vga_com_tile_module_n_178, B => vga_com_tile_module_n_265, C => vga_com_tile_module_n_52, ZN => vga_com_tile_module_n_545);
  vga_com_tile_module_g48177 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_347, A2 => vga_com_tile_module_n_92, B => vga_com_tile_module_n_10, Z => vga_com_tile_module_n_544);
  vga_com_tile_module_g48178 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_220, A2 => FE_OFN3_vga_com_row_1, B => vga_com_tile_module_n_442, ZN => vga_com_tile_module_n_543);
  vga_com_tile_module_g48179 : AOI211XD0BWP7T port map(A1 => vga_com_tile_module_n_18, A2 => vga_com_tile_module_n_15, B => vga_com_tile_module_n_289, C => vga_com_tile_module_n_180, ZN => vga_com_tile_module_n_542);
  vga_com_tile_module_g48180 : IOA21D1BWP7T port map(A1 => vga_com_tile_module_n_275, A2 => vga_com_tile_module_n_27, B => vga_com_tile_module_n_369, ZN => vga_com_tile_module_n_541);
  vga_com_tile_module_g48181 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_280, A2 => vga_com_tile_module_n_185, B1 => vga_com_tile_module_n_313, B2 => vga_com_tile_module_n_117, ZN => vga_com_tile_module_n_540);
  vga_com_tile_module_g48182 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_312, A2 => vga_com_tile_module_n_19, B1 => vga_com_tile_module_n_27, B2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_539);
  vga_com_tile_module_g48183 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_161, A2 => vga_com_tile_module_n_20, B => vga_com_tile_module_n_37, C => vga_com_tile_module_n_178, ZN => vga_com_tile_module_n_538);
  vga_com_tile_module_g48184 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_260, A2 => FE_OFN4_vga_com_row_2, B => vga_com_tile_module_n_16, ZN => vga_com_tile_module_n_537);
  vga_com_tile_module_g48185 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_133, A2 => vga_com_tile_module_n_368, B1 => vga_com_tile_module_n_166, B2 => vga_com_tile_module_n_251, ZN => vga_com_tile_module_n_536);
  vga_com_tile_module_g48186 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_316, A2 => vga_com_tile_module_n_28, B => vga_com_tile_module_n_187, ZN => vga_com_tile_module_n_535);
  vga_com_tile_module_g48187 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_314, A2 => vga_com_tile_module_n_208, B => vga_com_tile_module_n_126, Z => vga_com_tile_module_n_534);
  vga_com_tile_module_g48188 : IAO21D0BWP7T port map(A1 => vga_com_tile_module_n_319, A2 => vga_com_tile_module_n_275, B => vga_com_tile_module_n_122, ZN => vga_com_tile_module_n_533);
  vga_com_tile_module_g48189 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_340, A2 => vga_com_tile_module_n_65, B => vga_com_tile_module_n_26, ZN => vga_com_tile_module_n_532);
  vga_com_tile_module_g48190 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_256, A2 => vga_com_tile_module_n_27, B1 => vga_com_tile_module_n_183, B2 => vga_com_tile_module_n_106, ZN => vga_com_tile_module_n_531);
  vga_com_tile_module_g48191 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_471, A2 => vga_com_tile_module_n_22, ZN => vga_com_tile_module_n_530);
  vga_com_tile_module_g48192 : CKAN2D1BWP7T port map(A1 => vga_com_tile_module_n_444, A2 => vga_com_tile_module_n_29, Z => vga_com_tile_module_n_585);
  vga_com_tile_module_g48193 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_424, A2 => vga_com_tile_module_n_74, ZN => vga_com_tile_module_n_584);
  vga_com_tile_module_g48194 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_430, A2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_583);
  vga_com_tile_module_g48195 : AN2D0BWP7T port map(A1 => vga_com_tile_module_n_435, A2 => vga_com_tile_module_n_10, Z => vga_com_tile_module_n_582);
  vga_com_tile_module_g48196 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_427, A2 => vga_com_tile_module_n_432, ZN => vga_com_tile_module_n_581);
  vga_com_tile_module_g48197 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_367, A2 => vga_com_tile_module_n_9, B => vga_com_tile_module_n_413, Z => vga_com_tile_module_n_580);
  vga_com_tile_module_g48198 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_116, A2 => FE_OFN1_vga_com_row_0, B1 => vga_com_tile_module_n_8, B2 => vga_com_tile_module_n_47, C => vga_com_tile_module_n_175, ZN => vga_com_tile_module_n_579);
  vga_com_tile_module_g48199 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_428, A2 => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_529);
  vga_com_tile_module_g48200 : INR3D0BWP7T port map(A1 => vga_com_tile_module_n_363, B1 => FE_OFN3_vga_com_row_1, B2 => vga_com_tile_module_n_132, ZN => vga_com_tile_module_n_578);
  vga_com_tile_module_g48201 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_424, A2 => vga_com_tile_module_n_431, ZN => vga_com_tile_module_n_577);
  vga_com_tile_module_g48202 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_316, A2 => vga_com_tile_module_n_31, B => vga_com_tile_module_n_461, ZN => vga_com_tile_module_n_576);
  vga_com_tile_module_g48203 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_359, A2 => vga_com_tile_module_n_17, B1 => vga_com_tile_module_n_106, B2 => vga_com_tile_module_n_116, ZN => vga_com_tile_module_n_575);
  vga_com_tile_module_g48204 : OAI221D0BWP7T port map(A1 => vga_com_tile_module_n_211, A2 => vga_com_timer1(5), B1 => vga_com_tile_module_n_14, B2 => vga_com_tile_module_n_66, C => vga_com_tile_module_n_234, ZN => vga_com_tile_module_n_574);
  vga_com_tile_module_g48205 : AOI211D1BWP7T port map(A1 => vga_com_tile_module_n_51, A2 => vga_com_tile_module_n_9, B => vga_com_tile_module_n_306, C => vga_com_tile_module_n_65, ZN => vga_com_tile_module_n_573);
  vga_com_tile_module_g48206 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_315, A2 => vga_com_tile_module_n_295, B => vga_com_tile_module_n_391, ZN => vga_com_tile_module_n_572);
  vga_com_tile_module_g48207 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_424, A2 => vga_com_tile_module_n_192, ZN => vga_com_tile_module_n_571);
  vga_com_tile_module_g48208 : AOI221D1BWP7T port map(A1 => vga_com_tile_module_n_210, A2 => vga_com_timer1(5), B1 => vga_com_tile_module_n_67, B2 => vga_com_tile_module_n_14, C => vga_com_tile_module_n_233, ZN => vga_com_tile_module_n_569);
  vga_com_tile_module_g48209 : AOI31D1BWP7T port map(A1 => vga_com_tile_module_n_7, A2 => vga_com_bg_select(2), A3 => vga_com_bg_select(1), B => vga_com_tile_module_n_100, ZN => vga_com_tile_module_n_568);
  vga_com_tile_module_g48210 : INVD0BWP7T port map(I => vga_com_tile_module_n_525, ZN => vga_com_tile_module_n_526);
  vga_com_tile_module_g48211 : OA222D0BWP7T port map(A1 => vga_com_tile_module_n_228, A2 => vga_com_tile_module_n_30, B1 => vga_com_tile_module_n_21, B2 => vga_com_tile_module_n_201, C1 => vga_com_tile_module_n_10, C2 => vga_com_tile_module_n_246, Z => vga_com_tile_module_n_524);
  vga_com_tile_module_g48212 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_332, A2 => vga_com_tile_module_n_103, B1 => vga_com_tile_module_n_187, B2 => vga_com_tile_module_n_211, C1 => vga_com_tile_module_n_66, C2 => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_523);
  vga_com_tile_module_g48213 : AOI222D0BWP7T port map(A1 => vga_com_tile_module_n_314, A2 => vga_com_tile_module_n_113, B1 => vga_com_tile_module_n_176, B2 => vga_com_tile_module_n_185, C1 => vga_com_tile_module_n_182, C2 => vga_com_tile_module_n_103, ZN => vga_com_tile_module_n_522);
  vga_com_tile_module_g48214 : AOI32D1BWP7T port map(A1 => vga_com_tile_module_n_113, A2 => vga_com_tile_module_n_205, A3 => vga_com_tile_module_n_47, B1 => vga_com_tile_module_n_355, B2 => vga_com_tile_module_n_185, ZN => vga_com_tile_module_n_521);
  vga_com_tile_module_g48215 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_238, A2 => vga_com_tile_module_n_24, B1 => vga_com_tile_module_n_266, B2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_520);
  vga_com_tile_module_g48216 : OA22D0BWP7T port map(A1 => vga_com_tile_module_n_339, A2 => vga_com_tile_module_n_184, B1 => vga_com_tile_module_n_72, B2 => vga_com_tile_module_n_61, Z => vga_com_tile_module_n_519);
  vga_com_tile_module_g48217 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_351, A2 => vga_com_tile_module_n_231, B1 => vga_com_tile_module_n_162, B2 => vga_com_tile_module_n_46, ZN => vga_com_tile_module_n_518);
  vga_com_tile_module_g48218 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_346, A2 => vga_com_tile_module_n_30, B1 => vga_com_tile_module_n_339, B2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_517);
  vga_com_tile_module_g48219 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_276, A2 => vga_com_tile_module_n_10, B1 => vga_com_tile_module_n_74, B2 => vga_com_tile_module_n_21, ZN => vga_com_tile_module_n_516);
  vga_com_tile_module_g48220 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_148, A2 => vga_com_tile_module_n_278, B1 => vga_com_tile_module_n_202, B2 => vga_com_tile_module_n_245, ZN => vga_com_tile_module_n_515);
  vga_com_tile_module_g48221 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_145, A2 => vga_com_tile_module_n_235, B1 => vga_com_tile_module_n_326, B2 => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_514);
  vga_com_tile_module_g48222 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_281, A2 => vga_com_tile_module_n_334, B1 => vga_com_tile_module_n_344, B2 => vga_com_tile_module_n_193, ZN => vga_com_tile_module_n_513);
  vga_com_tile_module_g48223 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_20, A2 => vga_com_tile_module_n_85, B1 => vga_com_tile_module_n_337, B2 => vga_com_tile_module_n_30, ZN => vga_com_tile_module_n_512);
  vga_com_tile_module_g48224 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_286, A2 => vga_com_tile_module_n_27, B1 => vga_com_tile_module_n_28, B2 => vga_com_tile_module_n_64, ZN => vga_com_tile_module_n_511);
  vga_com_tile_module_g48225 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_353, A2 => vga_com_tile_module_n_185, B1 => vga_com_tile_module_n_109, B2 => vga_com_tile_module_n_75, ZN => vga_com_tile_module_n_510);
  vga_com_tile_module_g48226 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_154, A2 => vga_com_tile_module_n_361, B1 => vga_com_tile_module_n_147, B2 => vga_com_tile_module_n_66, ZN => vga_com_tile_module_n_509);
  vga_com_tile_module_g48227 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_316, A2 => vga_com_tile_module_n_25, B1 => vga_com_tile_module_n_258, B2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_508);
  vga_com_tile_module_g48228 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_265, A2 => vga_com_tile_module_n_185, B1 => vga_com_tile_module_n_361, B2 => vga_com_tile_module_n_111, ZN => vga_com_tile_module_n_507);
  vga_com_tile_module_g48229 : OA22D0BWP7T port map(A1 => vga_com_tile_module_n_288, A2 => vga_com_tile_module_n_18, B1 => vga_com_tile_module_n_29, B2 => vga_com_tile_module_n_350, Z => vga_com_tile_module_n_506);
  vga_com_tile_module_g48230 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_292, A2 => vga_com_tile_module_n_59, B1 => vga_com_tile_module_n_150, B2 => vga_com_tile_module_n_226, ZN => vga_com_tile_module_n_505);
  vga_com_tile_module_g48231 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_272, A2 => vga_com_tile_module_n_29, B1 => vga_com_tile_module_n_333, B2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_504);
  vga_com_tile_module_g48232 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_320, A2 => vga_com_tile_module_n_8, B1 => vga_com_tile_module_n_181, B2 => vga_com_tile_module_n_24, ZN => vga_com_tile_module_n_503);
  vga_com_tile_module_g48233 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_342, A2 => vga_com_tile_module_n_9, B1 => vga_com_tile_module_n_204, B2 => vga_com_tile_module_n_29, ZN => vga_com_tile_module_n_502);
  vga_com_tile_module_g48234 : AO22D0BWP7T port map(A1 => vga_com_tile_module_n_279, A2 => vga_com_tile_module_n_19, B1 => vga_com_tile_module_n_348, B2 => vga_com_tile_module_n_182, Z => vga_com_tile_module_n_501);
  vga_com_tile_module_g48235 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_281, A2 => vga_com_tile_module_n_23, B1 => vga_com_tile_module_n_213, B2 => vga_com_tile_module_n_21, ZN => vga_com_tile_module_n_500);
  vga_com_tile_module_g48236 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_127, A2 => vga_com_tile_module_n_364, B1 => vga_com_tile_module_n_150, B2 => vga_com_tile_module_n_353, ZN => vga_com_tile_module_n_499);
  vga_com_tile_module_g48237 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_347, A2 => vga_com_tile_module_n_16, B1 => vga_com_tile_module_n_144, B2 => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_498);
  vga_com_tile_module_g48238 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_319, A2 => vga_com_tile_module_n_9, B1 => vga_com_tile_module_n_365, B2 => vga_com_tile_module_n_26, ZN => vga_com_tile_module_n_497);
  vga_com_tile_module_g48239 : OA22D0BWP7T port map(A1 => vga_com_tile_module_n_279, A2 => vga_com_tile_module_n_110, B1 => vga_com_tile_module_n_207, B2 => vga_com_tile_module_n_112, Z => vga_com_tile_module_n_496);
  vga_com_tile_module_g48240 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_133, A2 => vga_com_tile_module_n_336, B1 => vga_com_tile_module_n_152, B2 => vga_com_tile_module_n_266, ZN => vga_com_tile_module_n_495);
  vga_com_tile_module_g48241 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_143, A2 => vga_com_tile_module_n_358, B1 => vga_com_tile_module_n_335, B2 => vga_com_tile_module_n_66, ZN => vga_com_tile_module_n_494);
  vga_com_tile_module_g48242 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_258, A2 => vga_com_tile_module_n_30, B1 => vga_com_tile_module_n_316, B2 => vga_com_tile_module_n_24, ZN => vga_com_tile_module_n_493);
  vga_com_tile_module_g48243 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_32, A2 => vga_com_tile_module_n_64, B1 => vga_com_tile_module_n_34, B2 => vga_com_tile_module_n_272, ZN => vga_com_tile_module_n_492);
  vga_com_tile_module_g48244 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_126, A2 => vga_com_tile_module_n_318, B1 => vga_com_tile_module_n_124, B2 => vga_com_tile_module_n_161, ZN => vga_com_tile_module_n_491);
  vga_com_tile_module_g48245 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_347, A2 => vga_com_tile_module_n_18, B1 => vga_com_tile_module_n_314, B2 => vga_com_tile_module_n_294, ZN => vga_com_tile_module_n_490);
  vga_com_tile_module_g48246 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_332, A2 => vga_com_tile_module_n_187, B1 => vga_com_tile_module_n_207, B2 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_489);
  vga_com_tile_module_g48247 : OA22D0BWP7T port map(A1 => vga_com_tile_module_n_327, A2 => vga_com_tile_module_n_143, B1 => vga_com_tile_module_n_183, B2 => vga_com_tile_module_n_150, Z => vga_com_tile_module_n_488);
  vga_com_tile_module_g48248 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_338, A2 => vga_com_tile_module_n_18, B1 => vga_com_tile_module_n_132, B2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_487);
  vga_com_tile_module_g48249 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_288, A2 => vga_com_tile_module_n_160, B1 => vga_com_tile_module_n_162, B2 => vga_com_tile_module_n_325, ZN => vga_com_tile_module_n_486);
  vga_com_tile_module_g48250 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_336, A2 => vga_com_tile_module_n_10, B1 => vga_com_tile_module_n_182, B2 => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_485);
  vga_com_tile_module_g48251 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_271, A2 => vga_com_tile_module_n_203, B1 => vga_com_tile_module_n_131, B2 => vga_com_tile_module_n_67, ZN => vga_com_tile_module_n_484);
  vga_com_tile_module_g48252 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_279, A2 => vga_com_tile_module_n_129, B1 => vga_com_tile_module_n_292, B2 => vga_com_tile_module_n_325, ZN => vga_com_tile_module_n_483);
  vga_com_tile_module_g48253 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_307, A2 => vga_com_tile_module_n_180, B1 => vga_com_tile_module_n_186, B2 => vga_com_tile_module_n_140, ZN => vga_com_tile_module_n_482);
  vga_com_tile_module_g48254 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_111, A2 => vga_com_tile_module_n_41, B1 => vga_com_tile_module_n_329, B2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_481);
  vga_com_tile_module_g48255 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_280, A2 => vga_com_tile_module_n_124, B1 => vga_com_tile_module_n_36, B2 => vga_com_tile_module_n_64, ZN => vga_com_tile_module_n_480);
  vga_com_tile_module_g48256 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_147, A2 => vga_com_tile_module_n_281, B1 => vga_com_tile_module_n_155, B2 => vga_com_tile_module_n_265, ZN => vga_com_tile_module_n_479);
  vga_com_tile_module_g48257 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_131, A2 => vga_com_tile_module_n_191, B1 => vga_com_tile_module_n_153, B2 => vga_com_tile_module_n_281, ZN => vga_com_tile_module_n_478);
  vga_com_tile_module_g48258 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_141, A2 => vga_com_tile_module_n_120, B1 => vga_com_tile_module_n_338, B2 => vga_com_tile_module_n_123, ZN => vga_com_tile_module_n_477);
  vga_com_tile_module_g48259 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_293, A2 => vga_com_tile_module_n_278, B1 => vga_com_tile_module_n_180, B2 => vga_com_tile_module_n_117, ZN => vga_com_tile_module_n_476);
  vga_com_tile_module_g48260 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_262, A2 => vga_com_tile_module_n_185, B1 => vga_com_tile_module_n_196, B2 => vga_com_tile_module_n_106, ZN => vga_com_tile_module_n_475);
  vga_com_tile_module_g48261 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_264, A2 => vga_com_tile_module_n_50, B1 => vga_com_tile_module_n_359, B2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_474);
  vga_com_tile_module_g48262 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_202, A2 => vga_com_tile_module_n_121, B1 => vga_com_tile_module_n_329, B2 => vga_com_tile_module_n_16, ZN => vga_com_tile_module_n_473);
  vga_com_tile_module_g48263 : MOAI22D0BWP7T port map(A1 => vga_com_tile_module_n_273, A2 => vga_com_tile_module_n_29, B1 => vga_com_tile_module_n_319, B2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_528);
  vga_com_tile_module_g48265 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_366, A2 => vga_com_tile_module_n_8, B1 => vga_com_tile_module_n_358, B2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_525);
  vga_com_tile_module_g48267 : INVD0BWP7T port map(I => vga_com_tile_module_n_451, ZN => vga_com_tile_module_n_452);
  vga_com_tile_module_g48268 : INVD0BWP7T port map(I => vga_com_tile_module_n_443, ZN => vga_com_tile_module_n_442);
  vga_com_tile_module_g48269 : INVD0BWP7T port map(I => vga_com_tile_module_n_441, ZN => vga_com_tile_module_n_440);
  vga_com_tile_module_g48270 : INVD0BWP7T port map(I => vga_com_tile_module_n_438, ZN => vga_com_tile_module_n_439);
  vga_com_tile_module_g48271 : INVD1BWP7T port map(I => vga_com_tile_module_n_433, ZN => vga_com_tile_module_n_434);
  vga_com_tile_module_g48272 : INVD0BWP7T port map(I => vga_com_tile_module_n_432, ZN => vga_com_tile_module_n_431);
  vga_com_tile_module_g48273 : INVD0BWP7T port map(I => vga_com_tile_module_n_430, ZN => vga_com_tile_module_n_429);
  vga_com_tile_module_g48274 : INVD0BWP7T port map(I => vga_com_tile_module_n_427, ZN => vga_com_tile_module_n_426);
  vga_com_tile_module_g48275 : INVD1BWP7T port map(I => vga_com_tile_module_n_425, ZN => vga_com_tile_module_n_424);
  vga_com_tile_module_g48276 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_272, A2 => vga_com_tile_module_n_104, ZN => vga_com_tile_module_n_423);
  vga_com_tile_module_g48277 : AN2D0BWP7T port map(A1 => vga_com_tile_module_n_367, A2 => vga_com_tile_module_n_121, Z => vga_com_tile_module_n_422);
  vga_com_tile_module_g48278 : CKND2D0BWP7T port map(A1 => vga_com_tile_module_n_351, A2 => vga_com_tile_module_n_193, ZN => vga_com_tile_module_n_421);
  vga_com_tile_module_g48279 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_326, A2 => vga_com_tile_module_n_140, ZN => vga_com_tile_module_n_420);
  vga_com_tile_module_g48280 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_277, A2 => vga_com_tile_module_n_273, ZN => vga_com_tile_module_n_472);
  vga_com_tile_module_g48281 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_259, A2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_471);
  vga_com_tile_module_g48282 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_361, A2 => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_419);
  vga_com_tile_module_g48283 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_362, A2 => vga_com_tile_module_n_18, Z => vga_com_tile_module_n_470);
  vga_com_tile_module_g48284 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_360, B1 => vga_com_tile_module_n_36, ZN => vga_com_tile_module_n_469);
  vga_com_tile_module_g48285 : AN2D0BWP7T port map(A1 => vga_com_tile_module_n_330, A2 => vga_com_tile_module_n_22, Z => vga_com_tile_module_n_468);
  vga_com_tile_module_g48286 : INR2D1BWP7T port map(A1 => vga_com_tile_module_n_330, B1 => vga_com_tile_module_n_178, ZN => vga_com_tile_module_n_467);
  vga_com_tile_module_g48287 : AN2D1BWP7T port map(A1 => vga_com_tile_module_n_273, A2 => vga_com_tile_module_n_121, Z => vga_com_tile_module_n_466);
  vga_com_tile_module_g48288 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_262, A2 => vga_com_tile_module_n_16, ZN => vga_com_tile_module_n_465);
  vga_com_tile_module_g48289 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_283, B1 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_464);
  vga_com_tile_module_g48290 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_340, A2 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_463);
  vga_com_tile_module_g48291 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_327, A2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_462);
  vga_com_tile_module_g48292 : AN2D0BWP7T port map(A1 => vga_com_tile_module_n_275, A2 => FE_OFN3_vga_com_row_1, Z => vga_com_tile_module_n_461);
  vga_com_tile_module_g48293 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_304, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_460);
  vga_com_tile_module_g48294 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_103, A2 => vga_com_tile_module_n_325, ZN => vga_com_tile_module_n_459);
  vga_com_tile_module_g48295 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_266, A2 => vga_com_tile_module_n_16, Z => vga_com_tile_module_n_458);
  vga_com_tile_module_g48296 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_259, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_457);
  vga_com_tile_module_g48297 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_189, A2 => vga_com_tile_module_n_276, ZN => vga_com_tile_module_n_456);
  vga_com_tile_module_g48298 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_260, A2 => vga_com_tile_module_n_144, ZN => vga_com_tile_module_n_455);
  vga_com_tile_module_g48299 : IND2D0BWP7T port map(A1 => vga_com_tile_module_n_144, B1 => vga_com_tile_module_n_273, ZN => vga_com_tile_module_n_454);
  vga_com_tile_module_g48300 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_304, A2 => vga_com_tile_module_n_32, ZN => vga_com_tile_module_n_453);
  vga_com_tile_module_g48301 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_322, A2 => vga_com_tile_module_n_191, ZN => vga_com_tile_module_n_451);
  vga_com_tile_module_g48302 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_322, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_450);
  vga_com_tile_module_g48303 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_315, A2 => vga_com_tile_module_n_113, ZN => vga_com_tile_module_n_449);
  vga_com_tile_module_g48304 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_280, A2 => vga_com_tile_module_n_204, Z => vga_com_tile_module_n_448);
  vga_com_tile_module_g48305 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_336, A2 => vga_com_tile_module_n_51, ZN => vga_com_tile_module_n_447);
  vga_com_tile_module_g48306 : INR2XD0BWP7T port map(A1 => vga_com_tile_module_n_207, B1 => vga_com_tile_module_n_350, ZN => vga_com_tile_module_n_446);
  vga_com_tile_module_g48307 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_315, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_445);
  vga_com_tile_module_g48308 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_261, A2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_444);
  vga_com_tile_module_g48309 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_289, B1 => vga_com_tile_module_n_156, ZN => vga_com_tile_module_n_443);
  vga_com_tile_module_g48310 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_262, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_441);
  vga_com_tile_module_g48311 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_329, A2 => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_438);
  vga_com_tile_module_g48312 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_336, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_437);
  vga_com_tile_module_g48314 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_293, A2 => vga_com_tile_module_n_263, ZN => vga_com_tile_module_n_436);
  vga_com_tile_module_g48315 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_182, A2 => vga_com_tile_module_n_323, ZN => vga_com_tile_module_n_435);
  vga_com_tile_module_g48316 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_326, A2 => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_433);
  vga_com_tile_module_g48317 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_362, A2 => vga_com_tile_module_n_179, ZN => vga_com_tile_module_n_432);
  vga_com_tile_module_g48318 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_336, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_430);
  vga_com_tile_module_g48319 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_324, A2 => vga_com_tile_module_n_77, ZN => vga_com_tile_module_n_428);
  vga_com_tile_module_g48320 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_172, A2 => vga_com_bg_select(0), ZN => vga_com_tile_module_n_427);
  vga_com_tile_module_g48321 : NR3D1BWP7T port map(A1 => vga_com_bg_select(0), A2 => vga_com_bg_select(2), A3 => vga_com_bg_select(1), ZN => vga_com_tile_module_n_425);
  vga_com_tile_module_g48322 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_108, A2 => vga_com_tile_module_n_127, A3 => vga_com_tile_module_n_139, ZN => vga_com_tile_module_n_411);
  vga_com_tile_module_g48323 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_164, A2 => vga_com_tile_module_n_23, B1 => vga_com_tile_module_n_78, B2 => vga_com_tile_module_n_21, ZN => vga_com_tile_module_n_410);
  vga_com_tile_module_g48324 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_220, A2 => vga_com_tile_module_n_9, B => vga_com_tile_module_n_26, ZN => vga_com_tile_module_n_409);
  vga_com_tile_module_g48325 : IAO21D0BWP7T port map(A1 => vga_com_tile_module_n_223, A2 => vga_com_tile_module_n_8, B => vga_com_tile_module_n_289, ZN => vga_com_tile_module_n_408);
  vga_com_tile_module_g48326 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_103, A2 => vga_com_tile_module_n_62, B1 => vga_com_tile_module_n_209, B2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_407);
  vga_com_tile_module_g48327 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_142, A2 => vga_com_tile_module_n_176, B1 => vga_com_tile_module_n_143, B2 => vga_com_tile_module_n_72, ZN => vga_com_tile_module_n_406);
  vga_com_tile_module_g48328 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_121, A2 => vga_com_tile_module_n_19, B1 => vga_com_tile_module_n_57, B2 => vga_com_tile_module_n_88, ZN => vga_com_tile_module_n_405);
  vga_com_tile_module_g48329 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_195, A2 => vga_com_tile_module_n_9, B => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_404);
  vga_com_tile_module_g48330 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_187, A2 => vga_com_tile_module_n_19, B => vga_com_tile_module_n_81, ZN => vga_com_tile_module_n_403);
  vga_com_tile_module_g48331 : AO211D0BWP7T port map(A1 => vga_com_tile_module_n_23, A2 => vga_com_tile_module_n_21, B => vga_com_tile_module_n_236, C => vga_com_tile_module_n_198, Z => vga_com_tile_module_n_402);
  vga_com_tile_module_g48332 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_120, A2 => FE_OFN3_vga_com_row_1, B1 => vga_com_tile_module_n_243, B2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_401);
  vga_com_tile_module_g48333 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_225, A2 => vga_com_tile_module_n_21, B1 => vga_com_tile_module_n_66, B2 => vga_com_tile_module_n_30, ZN => vga_com_tile_module_n_400);
  vga_com_tile_module_g48334 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_183, A2 => vga_com_tile_module_n_76, B => vga_com_tile_module_n_103, ZN => vga_com_tile_module_n_399);
  vga_com_tile_module_g48335 : NR3D0BWP7T port map(A1 => vga_com_tile_module_n_196, A2 => vga_com_tile_module_n_104, A3 => vga_com_tile_module_n_79, ZN => vga_com_tile_module_n_398);
  vga_com_tile_module_g48336 : MAOI22D0BWP7T port map(A1 => vga_com_tile_module_n_65, A2 => vga_com_tile_module_n_57, B1 => vga_com_tile_module_n_213, B2 => vga_com_tile_module_n_53, ZN => vga_com_tile_module_n_397);
  vga_com_tile_module_g48337 : ND3D0BWP7T port map(A1 => vga_com_tile_module_n_127, A2 => vga_com_tile_module_n_204, A3 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_396);
  vga_com_tile_module_g48338 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_179, A2 => FE_OFN4_vga_com_row_2, B => vga_com_tile_module_n_29, ZN => vga_com_tile_module_n_395);
  vga_com_tile_module_g48339 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_190, A2 => vga_com_tile_module_n_80, B => vga_com_tile_module_n_130, ZN => vga_com_tile_module_n_394);
  vga_com_tile_module_g48340 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_215, A2 => vga_com_tile_module_n_29, B => vga_com_tile_module_n_104, ZN => vga_com_tile_module_n_393);
  vga_com_tile_module_g48341 : IOA21D1BWP7T port map(A1 => vga_com_tile_module_n_140, A2 => vga_com_tile_module_n_17, B => vga_com_tile_module_n_110, ZN => vga_com_tile_module_n_392);
  vga_com_tile_module_g48342 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_118, A2 => vga_com_tile_module_n_104, B => vga_com_tile_module_n_73, ZN => vga_com_tile_module_n_391);
  vga_com_tile_module_g48343 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_219, A2 => vga_com_tile_module_n_16, B => vga_com_tile_module_n_266, ZN => vga_com_tile_module_n_390);
  vga_com_tile_module_g48344 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_181, A2 => vga_com_tile_module_n_30, B => vga_com_tile_module_n_330, Z => vga_com_tile_module_n_389);
  vga_com_tile_module_g48345 : IOA21D0BWP7T port map(A1 => vga_com_tile_module_n_222, A2 => vga_com_tile_module_n_12, B => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_388);
  vga_com_tile_module_g48346 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_196, A2 => vga_com_tile_module_n_8, B => vga_com_tile_module_n_239, ZN => vga_com_tile_module_n_387);
  vga_com_tile_module_g48347 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_139, A2 => vga_com_tile_module_n_124, B => vga_com_tile_module_n_194, ZN => vga_com_tile_module_n_386);
  vga_com_tile_module_g48348 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_138, A2 => vga_com_tile_module_n_129, B => vga_com_tile_module_n_46, ZN => vga_com_tile_module_n_385);
  vga_com_tile_module_g48349 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_182, A2 => vga_com_tile_module_n_181, B => vga_com_tile_module_n_114, ZN => vga_com_tile_module_n_384);
  vga_com_tile_module_g48350 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_206, A2 => vga_com_tile_module_n_72, B => vga_com_tile_module_n_22, Z => vga_com_tile_module_n_383);
  vga_com_tile_module_g48351 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_218, A2 => FE_OFN3_vga_com_row_1, B => vga_com_tile_module_n_22, ZN => vga_com_tile_module_n_382);
  vga_com_tile_module_g48352 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_125, A2 => vga_com_tile_module_n_129, B => vga_com_tile_module_n_269, ZN => vga_com_tile_module_n_381);
  vga_com_tile_module_g48353 : IND3D0BWP7T port map(A1 => vga_com_tile_module_n_212, B1 => vga_com_tile_module_n_47, B2 => vga_com_tile_module_n_127, ZN => vga_com_tile_module_n_380);
  vga_com_tile_module_g48354 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_118, A2 => vga_com_tile_module_n_112, B => vga_com_tile_module_n_269, ZN => vga_com_tile_module_n_379);
  vga_com_tile_module_g48355 : MAOI22D0BWP7T port map(A1 => vga_com_column(2), A2 => vga_com_timer1(5), B1 => vga_com_tile_module_n_206, B2 => vga_com_timer1(5), ZN => vga_com_tile_module_n_378);
  vga_com_tile_module_g48356 : MAOI22D0BWP7T port map(A1 => vga_com_column(2), A2 => vga_com_tile_module_n_14, B1 => vga_com_tile_module_n_206, B2 => vga_com_tile_module_n_14, ZN => vga_com_tile_module_n_377);
  vga_com_tile_module_g48357 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_185, A2 => vga_com_tile_module_n_224, B1 => vga_com_tile_module_n_187, B2 => vga_com_tile_module_n_77, ZN => vga_com_tile_module_n_376);
  vga_com_tile_module_g48358 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_113, A2 => vga_com_tile_module_n_224, B1 => vga_com_tile_module_n_197, B2 => vga_com_tile_module_n_57, ZN => vga_com_tile_module_n_375);
  vga_com_tile_module_g48359 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_118, A2 => vga_com_column(1), B1 => vga_com_tile_module_n_41, B2 => vga_com_tile_module_n_53, ZN => vga_com_tile_module_n_374);
  vga_com_tile_module_g48360 : AOI22D0BWP7T port map(A1 => vga_com_tile_module_n_217, A2 => vga_com_tile_module_n_111, B1 => vga_com_tile_module_n_52, B2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_373);
  vga_com_tile_module_g48361 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_200, A2 => FE_OFN1_vga_com_row_0, B => vga_com_tile_module_n_91, ZN => vga_com_tile_module_n_418);
  vga_com_tile_module_g48362 : ND3D0BWP7T port map(A1 => vga_com_tile_module_n_123, A2 => vga_com_tile_module_n_216, A3 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_417);
  vga_com_tile_module_g48363 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_41, A2 => FE_OFN1_vga_com_row_0, B => vga_com_tile_module_n_274, ZN => vga_com_tile_module_n_416);
  vga_com_tile_module_g48364 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_196, A2 => FE_OFN1_vga_com_row_0, B => vga_com_tile_module_n_333, ZN => vga_com_tile_module_n_415);
  vga_com_tile_module_g48365 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_200, A2 => FE_OFN3_vga_com_row_1, B => vga_com_tile_module_n_21, ZN => vga_com_tile_module_n_414);
  vga_com_tile_module_g48366 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_73, A2 => FE_OFN4_vga_com_row_2, B => vga_com_tile_module_n_306, Z => vga_com_tile_module_n_413);
  vga_com_tile_module_g48367 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_199, A2 => FE_OFN1_vga_com_row_0, B => vga_com_tile_module_n_319, ZN => vga_com_tile_module_n_412);
  vga_com_tile_module_g48369 : INVD0BWP7T port map(I => vga_com_tile_module_n_345, ZN => vga_com_tile_module_n_346);
  vga_com_tile_module_g48370 : INVD0BWP7T port map(I => vga_com_tile_module_n_344, ZN => vga_com_tile_module_n_343);
  vga_com_tile_module_g48371 : INVD0BWP7T port map(I => vga_com_tile_module_n_335, ZN => vga_com_tile_module_n_334);
  vga_com_tile_module_g48372 : INVD0BWP7T port map(I => vga_com_tile_module_n_332, ZN => vga_com_tile_module_n_331);
  vga_com_tile_module_g48373 : INVD1BWP7T port map(I => vga_com_tile_module_n_328, ZN => vga_com_tile_module_n_327);
  vga_com_tile_module_g48374 : INVD1BWP7T port map(I => vga_com_tile_module_n_325, ZN => vga_com_tile_module_n_324);
  vga_com_tile_module_g48375 : INVD1BWP7T port map(I => vga_com_tile_module_n_323, ZN => vga_com_tile_module_n_322);
  vga_com_tile_module_g48376 : INVD1BWP7T port map(I => vga_com_tile_module_n_321, ZN => vga_com_tile_module_n_320);
  vga_com_tile_module_g48377 : INVD0BWP7T port map(I => vga_com_tile_module_n_319, ZN => vga_com_tile_module_n_318);
  vga_com_tile_module_g48378 : INVD1BWP7T port map(I => vga_com_tile_module_n_317, ZN => vga_com_tile_module_n_316);
  vga_com_tile_module_g48379 : INVD1BWP7T port map(I => vga_com_tile_module_n_315, ZN => vga_com_tile_module_n_314);
  vga_com_tile_module_g48380 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_207, A2 => vga_com_tile_module_n_85, ZN => vga_com_tile_module_n_313);
  vga_com_tile_module_g48381 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_195, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_312);
  vga_com_tile_module_g48382 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_183, A2 => vga_com_tile_module_n_218, ZN => vga_com_tile_module_n_311);
  vga_com_tile_module_g48383 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_132, A2 => vga_com_tile_module_n_88, ZN => vga_com_tile_module_n_310);
  vga_com_tile_module_g48384 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_220, B1 => vga_com_tile_module_n_203, ZN => vga_com_tile_module_n_372);
  vga_com_tile_module_g48385 : INR2XD0BWP7T port map(A1 => vga_com_tile_module_n_101, B1 => vga_com_tile_module_n_140, ZN => vga_com_tile_module_n_371);
  vga_com_tile_module_g48386 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_104, A2 => vga_com_column(1), ZN => vga_com_tile_module_n_370);
  vga_com_tile_module_g48387 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_103, A2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_369);
  vga_com_tile_module_g48388 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_140, A2 => vga_com_tile_module_n_204, Z => vga_com_tile_module_n_368);
  vga_com_tile_module_g48389 : CKND2D0BWP7T port map(A1 => vga_com_tile_module_n_183, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_367);
  vga_com_tile_module_g48390 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_228, A2 => vga_com_tile_module_n_178, ZN => vga_com_tile_module_n_366);
  vga_com_tile_module_g48391 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_192, A2 => vga_com_tile_module_n_59, ZN => vga_com_tile_module_n_365);
  vga_com_tile_module_g48392 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_207, A2 => vga_com_tile_module_n_8, Z => vga_com_tile_module_n_364);
  vga_com_tile_module_g48393 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_219, A2 => vga_com_tile_module_n_80, ZN => vga_com_tile_module_n_363);
  vga_com_tile_module_g48394 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_193, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_362);
  vga_com_tile_module_g48395 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_198, A2 => vga_com_tile_module_n_88, ZN => vga_com_tile_module_n_361);
  vga_com_tile_module_g48396 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_235, B1 => vga_com_tile_module_n_217, ZN => vga_com_tile_module_n_360);
  vga_com_tile_module_g48397 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_115, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_359);
  vga_com_tile_module_g48398 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_196, A2 => vga_com_tile_module_n_64, ZN => vga_com_tile_module_n_358);
  vga_com_tile_module_g48399 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_212, B1 => vga_com_tile_module_n_193, ZN => vga_com_tile_module_n_357);
  vga_com_tile_module_g48400 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_197, A2 => vga_com_tile_module_n_231, ZN => vga_com_tile_module_n_356);
  vga_com_tile_module_g48401 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_197, A2 => vga_com_tile_module_n_205, ZN => vga_com_tile_module_n_355);
  vga_com_tile_module_g48402 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_109, A2 => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_354);
  vga_com_tile_module_g48403 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_201, A2 => vga_com_tile_module_n_47, ZN => vga_com_tile_module_n_353);
  vga_com_tile_module_g48404 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_112, A2 => vga_com_tile_module_n_201, ZN => vga_com_tile_module_n_352);
  vga_com_tile_module_g48405 : NR2D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_112, ZN => vga_com_tile_module_n_351);
  vga_com_tile_module_g48406 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_115, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_350);
  vga_com_tile_module_g48407 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_178, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_349);
  vga_com_tile_module_g48408 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_222, A2 => vga_com_tile_module_n_26, ZN => vga_com_tile_module_n_348);
  vga_com_tile_module_g48409 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_193, A2 => vga_com_tile_module_n_67, ZN => vga_com_tile_module_n_347);
  vga_com_tile_module_g48410 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_225, A2 => vga_com_tile_module_n_41, ZN => vga_com_tile_module_n_345);
  vga_com_tile_module_g48411 : NR2D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_184, ZN => vga_com_tile_module_n_344);
  vga_com_tile_module_g48412 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_190, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_342);
  vga_com_tile_module_g48413 : INR2D1BWP7T port map(A1 => vga_com_tile_module_n_207, B1 => vga_com_tile_module_n_191, ZN => vga_com_tile_module_n_341);
  vga_com_tile_module_g48414 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_194, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_340);
  vga_com_tile_module_g48415 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_221, A2 => vga_com_tile_module_n_178, ZN => vga_com_tile_module_n_339);
  vga_com_tile_module_g48416 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_120, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_338);
  vga_com_tile_module_g48417 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_116, A2 => vga_com_tile_module_n_4, ZN => vga_com_tile_module_n_337);
  vga_com_tile_module_g48418 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_234, A2 => vga_com_tile_module_n_211, ZN => vga_com_tile_module_n_336);
  vga_com_tile_module_g48419 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_2, A2 => vga_com_tile_module_n_113, ZN => vga_com_tile_module_n_335);
  vga_com_tile_module_g48420 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_201, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_333);
  vga_com_tile_module_g48421 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_223, A2 => vga_com_tile_module_n_195, ZN => vga_com_tile_module_n_332);
  vga_com_tile_module_g48422 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_213, A2 => vga_com_tile_module_n_64, Z => vga_com_tile_module_n_330);
  vga_com_tile_module_g48423 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_191, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_329);
  vga_com_tile_module_g48424 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_206, A2 => vga_com_tile_module_n_11, ZN => vga_com_tile_module_n_328);
  vga_com_tile_module_g48425 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_178, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_326);
  vga_com_tile_module_g48426 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_116, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_325);
  vga_com_tile_module_g48427 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_116, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_323);
  vga_com_tile_module_g48428 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_205, A2 => vga_com_tile_module_n_224, ZN => vga_com_tile_module_n_321);
  vga_com_tile_module_g48429 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_181, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_319);
  vga_com_tile_module_g48430 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_116, A2 => vga_com_tile_module_n_81, ZN => vga_com_tile_module_n_317);
  vga_com_tile_module_g48431 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_218, A2 => vga_com_tile_module_n_213, ZN => vga_com_tile_module_n_315);
  vga_com_tile_module_g48432 : INVD0BWP7T port map(I => vga_com_tile_module_n_296, ZN => vga_com_tile_module_n_297);
  vga_com_tile_module_g48433 : INVD0BWP7T port map(I => vga_com_tile_module_n_286, ZN => vga_com_tile_module_n_287);
  vga_com_tile_module_g48434 : CKND1BWP7T port map(I => vga_com_tile_module_n_284, ZN => vga_com_tile_module_n_285);
  vga_com_tile_module_g48435 : INVD0BWP7T port map(I => vga_com_tile_module_n_275, ZN => vga_com_tile_module_n_274);
  vga_com_tile_module_g48436 : INVD0BWP7T port map(I => vga_com_tile_module_n_272, ZN => vga_com_tile_module_n_271);
  vga_com_tile_module_g48437 : INVD1BWP7T port map(I => vga_com_tile_module_n_270, ZN => vga_com_tile_module_n_269);
  vga_com_tile_module_g48438 : INVD0BWP7T port map(I => vga_com_tile_module_n_268, ZN => vga_com_tile_module_n_267);
  vga_com_tile_module_g48439 : INVD0BWP7T port map(I => vga_com_tile_module_n_265, ZN => vga_com_tile_module_n_264);
  vga_com_tile_module_g48440 : INVD1BWP7T port map(I => vga_com_tile_module_n_263, ZN => vga_com_tile_module_n_262);
  vga_com_tile_module_g48441 : INVD1BWP7T port map(I => vga_com_tile_module_n_261, ZN => vga_com_tile_module_n_260);
  vga_com_tile_module_g48442 : INVD0BWP7T port map(I => vga_com_tile_module_n_259, ZN => vga_com_tile_module_n_258);
  vga_com_tile_module_g48443 : AO21D0BWP7T port map(A1 => vga_com_tile_module_n_65, A2 => vga_com_tile_module_n_16, B => vga_com_tile_module_n_132, Z => vga_com_tile_module_n_257);
  vga_com_tile_module_g48444 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_219, A2 => vga_com_tile_module_n_62, Z => vga_com_tile_module_n_256);
  vga_com_tile_module_g48445 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_51, A2 => vga_com_tile_module_n_10, B => vga_com_tile_module_n_179, ZN => vga_com_tile_module_n_255);
  vga_com_tile_module_g48446 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_40, A2 => vga_com_tile_module_n_63, B => vga_com_tile_module_n_24, ZN => vga_com_tile_module_n_254);
  vga_com_tile_module_g48447 : AN3D0BWP7T port map(A1 => vga_com_tile_module_n_36, A2 => vga_com_tile_module_n_173, A3 => vga_com_tile_module_n_51, Z => vga_com_tile_module_n_253);
  vga_com_tile_module_g48448 : OAI22D0BWP7T port map(A1 => vga_com_tile_module_n_41, A2 => vga_com_tile_module_n_30, B1 => vga_com_tile_module_n_23, B2 => vga_com_tile_module_n_79, ZN => vga_com_tile_module_n_252);
  vga_com_tile_module_g48449 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_206, A2 => vga_com_tile_module_n_67, ZN => vga_com_tile_module_n_251);
  vga_com_tile_module_g48450 : AN2D0BWP7T port map(A1 => vga_com_tile_module_n_125, A2 => vga_com_tile_module_n_143, Z => vga_com_tile_module_n_250);
  vga_com_tile_module_g48451 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_22, A2 => vga_com_tile_module_n_74, B => vga_com_tile_module_n_36, ZN => vga_com_tile_module_n_249);
  vga_com_tile_module_g48452 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_181, A2 => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_248);
  vga_com_tile_module_g48453 : IND2D0BWP7T port map(A1 => vga_com_tile_module_n_212, B1 => vga_com_tile_module_n_39, ZN => vga_com_tile_module_n_309);
  vga_com_tile_module_g48454 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_21, A2 => vga_com_column(2), B => vga_com_tile_module_n_192, ZN => vga_com_tile_module_n_308);
  vga_com_tile_module_g48455 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_17, A2 => vga_com_tile_module_n_63, B => vga_com_tile_module_n_109, ZN => vga_com_tile_module_n_307);
  vga_com_tile_module_g48456 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_18, A2 => vga_com_tile_module_n_51, B => vga_com_tile_module_n_16, ZN => vga_com_tile_module_n_306);
  vga_com_tile_module_g48457 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_191, A2 => vga_com_tile_module_n_105, ZN => vga_com_tile_module_n_305);
  vga_com_tile_module_g48458 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_197, A2 => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_304);
  vga_com_tile_module_g48459 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_107, A2 => vga_com_tile_module_n_136, ZN => vga_com_tile_module_n_303);
  vga_com_tile_module_g48460 : CKND2D0BWP7T port map(A1 => vga_com_tile_module_n_106, A2 => vga_com_tile_module_n_116, ZN => vga_com_tile_module_n_247);
  vga_com_tile_module_g48461 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_106, A2 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_302);
  vga_com_tile_module_g48462 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_168, A2 => vga_com_tile_module_n_21, Z => vga_com_tile_module_n_301);
  vga_com_tile_module_g48463 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_84, A2 => vga_com_tile_module_n_8, B => vga_com_tile_module_n_239, ZN => vga_com_tile_module_n_300);
  vga_com_tile_module_g48464 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_121, A2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_299);
  vga_com_tile_module_g48465 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_216, A2 => vga_com_tile_module_n_20, ZN => vga_com_tile_module_n_298);
  vga_com_tile_module_g48466 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_91, A2 => vga_com_tile_module_n_12, B => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_296);
  vga_com_tile_module_g48467 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_114, A2 => vga_com_tile_module_n_112, ZN => vga_com_tile_module_n_295);
  vga_com_tile_module_g48468 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_186, A2 => vga_com_tile_module_n_26, ZN => vga_com_tile_module_n_294);
  vga_com_tile_module_g48469 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_105, A2 => vga_com_tile_module_n_110, ZN => vga_com_tile_module_n_293);
  vga_com_tile_module_g48470 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_189, A2 => vga_com_tile_module_n_122, ZN => vga_com_tile_module_n_292);
  vga_com_tile_module_g48471 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_110, A2 => vga_com_tile_module_n_179, ZN => vga_com_tile_module_n_291);
  vga_com_tile_module_g48472 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_206, A2 => vga_com_tile_module_n_73, ZN => vga_com_tile_module_n_290);
  vga_com_tile_module_g48473 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_198, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_289);
  vga_com_tile_module_g48474 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_115, A2 => vga_com_tile_module_n_47, ZN => vga_com_tile_module_n_288);
  vga_com_tile_module_g48475 : AOI21D0BWP7T port map(A1 => vga_com_tile_module_n_75, A2 => FE_OFN1_vga_com_row_0, B => vga_com_column(2), ZN => vga_com_tile_module_n_286);
  vga_com_tile_module_g48476 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_121, A2 => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_284);
  vga_com_tile_module_g48477 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_119, A2 => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_283);
  vga_com_tile_module_g48478 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_137, B1 => vga_com_tile_module_n_136, ZN => vga_com_tile_module_n_282);
  vga_com_tile_module_g48479 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_115, A2 => vga_com_tile_module_n_40, ZN => vga_com_tile_module_n_281);
  vga_com_tile_module_g48480 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_140, B1 => vga_com_tile_module_n_85, ZN => vga_com_tile_module_n_280);
  vga_com_tile_module_g48481 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_183, A2 => vga_com_tile_module_n_119, ZN => vga_com_tile_module_n_279);
  vga_com_tile_module_g48482 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_179, A2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_278);
  vga_com_tile_module_g48483 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_196, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_277);
  vga_com_tile_module_g48484 : AOI21D0BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_column(1), B => vga_com_tile_module_n_195, ZN => vga_com_tile_module_n_276);
  vga_com_tile_module_g48485 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_191, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_275);
  vga_com_tile_module_g48486 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_180, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_273);
  vga_com_tile_module_g48487 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_178, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_272);
  vga_com_tile_module_g48488 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_181, A2 => vga_com_tile_module_n_195, ZN => vga_com_tile_module_n_270);
  vga_com_tile_module_g48489 : XNR2D1BWP7T port map(A1 => vga_com_tile_module_n_100, A2 => vga_com_bg_select(2), ZN => vga_com_tile_module_n_268);
  vga_com_tile_module_g48490 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_194, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_266);
  vga_com_tile_module_g48491 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_115, A2 => vga_com_tile_module_n_85, ZN => vga_com_tile_module_n_265);
  vga_com_tile_module_g48492 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_181, A2 => vga_com_tile_module_n_179, ZN => vga_com_tile_module_n_263);
  vga_com_tile_module_g48493 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_179, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_261);
  vga_com_tile_module_g48494 : AOI21D2BWP7T port map(A1 => vga_com_tile_module_n_67, A2 => vga_com_tile_module_n_4, B => vga_com_tile_module_n_228, ZN => vga_com_tile_module_n_259);
  vga_com_tile_module_g48495 : INVD0BWP7T port map(I => vga_com_tile_module_n_234, ZN => vga_com_tile_module_n_233);
  vga_com_tile_module_g48496 : CKND1BWP7T port map(I => vga_com_tile_module_n_231, ZN => vga_com_tile_module_n_232);
  vga_com_tile_module_g48497 : INVD0BWP7T port map(I => vga_com_tile_module_n_229, ZN => vga_com_tile_module_n_230);
  vga_com_tile_module_g48498 : INVD0BWP7T port map(I => vga_com_tile_module_n_218, ZN => vga_com_tile_module_n_217);
  vga_com_tile_module_g48499 : CKND1BWP7T port map(I => vga_com_tile_module_n_216, ZN => vga_com_tile_module_n_215);
  vga_com_tile_module_g48500 : INVD0BWP7T port map(I => vga_com_tile_module_n_211, ZN => vga_com_tile_module_n_210);
  vga_com_tile_module_g48501 : INVD0BWP7T port map(I => vga_com_tile_module_n_209, ZN => vga_com_tile_module_n_208);
  vga_com_tile_module_g48502 : INVD1BWP7T port map(I => vga_com_tile_module_n_205, ZN => vga_com_tile_module_n_204);
  vga_com_tile_module_g48503 : INVD0BWP7T port map(I => vga_com_tile_module_n_203, ZN => vga_com_tile_module_n_202);
  vga_com_tile_module_g48504 : INVD1BWP7T port map(I => vga_com_tile_module_n_201, ZN => vga_com_tile_module_n_200);
  vga_com_tile_module_g48505 : INVD1BWP7T port map(I => vga_com_tile_module_n_199, ZN => vga_com_tile_module_n_198);
  vga_com_tile_module_g48506 : INVD1BWP7T port map(I => vga_com_tile_module_n_197, ZN => vga_com_tile_module_n_196);
  vga_com_tile_module_g48507 : INVD1BWP7T port map(I => vga_com_tile_module_n_195, ZN => vga_com_tile_module_n_194);
  vga_com_tile_module_g48508 : INVD1BWP7T port map(I => vga_com_tile_module_n_193, ZN => vga_com_tile_module_n_192);
  vga_com_tile_module_g48509 : INVD1BWP7T port map(I => vga_com_tile_module_n_191, ZN => vga_com_tile_module_n_190);
  vga_com_tile_module_g48510 : INVD1BWP7T port map(I => vga_com_tile_module_n_189, ZN => vga_com_tile_module_n_188);
  vga_com_tile_module_g48511 : INVD1BWP7T port map(I => vga_com_tile_module_n_187, ZN => vga_com_tile_module_n_186);
  vga_com_tile_module_g48512 : INVD1BWP7T port map(I => vga_com_tile_module_n_185, ZN => vga_com_tile_module_n_184);
  vga_com_tile_module_g48513 : INVD1BWP7T port map(I => vga_com_tile_module_n_183, ZN => vga_com_tile_module_n_182);
  vga_com_tile_module_g48514 : INVD1BWP7T port map(I => vga_com_tile_module_n_181, ZN => vga_com_tile_module_n_180);
  vga_com_tile_module_g48515 : INVD1BWP7T port map(I => vga_com_tile_module_n_179, ZN => vga_com_tile_module_n_178);
  vga_com_tile_module_g48516 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_tile_module_n_81, ZN => vga_com_tile_module_n_177);
  vga_com_tile_module_g48517 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_tile_module_n_91, ZN => vga_com_tile_module_n_246);
  vga_com_tile_module_g48518 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_40, A2 => vga_com_tile_module_n_12, ZN => vga_com_tile_module_n_245);
  vga_com_tile_module_g48519 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_75, A2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_244);
  vga_com_tile_module_g48520 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_75, A2 => vga_com_tile_module_n_40, ZN => vga_com_tile_module_n_243);
  vga_com_tile_module_g48521 : CKND2D0BWP7T port map(A1 => vga_com_tile_module_n_45, A2 => vga_com_tile_module_n_5, ZN => vga_com_tile_module_n_242);
  vga_com_tile_module_g48522 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_95, A2 => vga_com_tile_module_n_3, Z => vga_com_tile_module_n_241);
  vga_com_tile_module_g48523 : OR2D1BWP7T port map(A1 => vga_com_tile_module_n_98, A2 => vga_com_tile_module_n_93, Z => vga_com_tile_module_n_240);
  vga_com_tile_module_g48524 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_80, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_239);
  vga_com_tile_module_g48525 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_87, A2 => vga_com_column(1), ZN => vga_com_tile_module_n_238);
  vga_com_tile_module_g48526 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_54, A2 => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_237);
  vga_com_tile_module_g48527 : ND2D1BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_34, ZN => vga_com_tile_module_n_236);
  vga_com_tile_module_g48528 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_235);
  vga_com_tile_module_g48529 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_67, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_234);
  vga_com_tile_module_g48530 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_63, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_231);
  vga_com_tile_module_g48531 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_5, A2 => vga_com_tile_module_n_94, ZN => vga_com_tile_module_n_229);
  vga_com_tile_module_g48532 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_tile_module_n_4, ZN => vga_com_tile_module_n_228);
  vga_com_tile_module_g48533 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_49, A2 => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_227);
  vga_com_tile_module_g48534 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_84, A2 => vga_com_column(2), ZN => vga_com_tile_module_n_226);
  vga_com_tile_module_g48535 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_67, A2 => vga_com_tile_module_n_77, ZN => vga_com_tile_module_n_225);
  vga_com_tile_module_g48536 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_40, A2 => vga_com_column(1), ZN => vga_com_tile_module_n_224);
  vga_com_tile_module_g48537 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_72, A2 => vga_com_tile_module_n_81, ZN => vga_com_tile_module_n_223);
  vga_com_tile_module_g48538 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_21, A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_222);
  vga_com_tile_module_g48539 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_77, A2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_221);
  vga_com_tile_module_g48540 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_76, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_220);
  vga_com_tile_module_g48541 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_219);
  vga_com_tile_module_g48542 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_72, A2 => vga_com_tile_module_n_4, ZN => vga_com_tile_module_n_218);
  vga_com_tile_module_g48543 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_88, A2 => vga_com_tile_module_n_67, ZN => vga_com_tile_module_n_216);
  vga_com_tile_module_g48544 : ND2D1BWP7T port map(A1 => vga_com_tile_address(2), A2 => vga_com_tile_module_n_94, ZN => vga_com_tile_module_n_214);
  vga_com_tile_module_g48545 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_88, A2 => vga_com_tile_module_n_75, ZN => vga_com_tile_module_n_213);
  vga_com_tile_module_g48546 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_77, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_212);
  vga_com_tile_module_g48547 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_73, A2 => vga_com_tile_module_n_4, ZN => vga_com_tile_module_n_211);
  vga_com_tile_module_g48548 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_80, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_209);
  vga_com_tile_module_g48549 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_79, A2 => vga_com_column(2), ZN => vga_com_tile_module_n_207);
  vga_com_tile_module_g48550 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_75, A2 => vga_com_tile_module_n_77, ZN => vga_com_tile_module_n_206);
  vga_com_tile_module_g48551 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_205);
  vga_com_tile_module_g48552 : NR2D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_18, ZN => vga_com_tile_module_n_203);
  vga_com_tile_module_g48553 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_76, A2 => vga_com_tile_module_n_11, ZN => vga_com_tile_module_n_201);
  vga_com_tile_module_g48554 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_63, A2 => vga_com_tile_module_n_80, ZN => vga_com_tile_module_n_199);
  vga_com_tile_module_g48555 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_62, A2 => vga_com_tile_module_n_4, ZN => vga_com_tile_module_n_197);
  vga_com_tile_module_g48556 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_77, A2 => vga_com_tile_module_n_11, ZN => vga_com_tile_module_n_195);
  vga_com_tile_module_g48557 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_77, A2 => vga_com_column(2), ZN => vga_com_tile_module_n_193);
  vga_com_tile_module_g48558 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_67, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_191);
  vga_com_tile_module_g48559 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_34, A2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_189);
  vga_com_tile_module_g48560 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_23, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_187);
  vga_com_tile_module_g48561 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_21, A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_185);
  vga_com_tile_module_g48562 : NR2D1P5BWP7T port map(A1 => vga_com_tile_module_n_73, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_183);
  vga_com_tile_module_g48563 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_62, A2 => vga_com_column(0), ZN => vga_com_tile_module_n_181);
  vga_com_tile_module_g48564 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_tile_module_n_4, ZN => vga_com_tile_module_n_179);
  vga_com_tile_module_g48565 : INVD0BWP7T port map(I => vga_com_tile_module_n_165, ZN => vga_com_tile_module_n_166);
  vga_com_tile_module_g48566 : CKND1BWP7T port map(I => vga_com_tile_module_n_163, ZN => vga_com_tile_module_n_164);
  vga_com_tile_module_g48567 : INVD0BWP7T port map(I => vga_com_tile_module_n_158, ZN => vga_com_tile_module_n_159);
  vga_com_tile_module_g48568 : INVD0BWP7T port map(I => vga_com_tile_module_n_155, ZN => vga_com_tile_module_n_154);
  vga_com_tile_module_g48569 : INVD0BWP7T port map(I => vga_com_tile_module_n_152, ZN => vga_com_tile_module_n_151);
  vga_com_tile_module_g48570 : INVD0BWP7T port map(I => vga_com_tile_module_n_149, ZN => vga_com_tile_module_n_148);
  vga_com_tile_module_g48571 : CKND1BWP7T port map(I => vga_com_tile_module_n_146, ZN => vga_com_tile_module_n_145);
  vga_com_tile_module_g48572 : INVD0BWP7T port map(I => vga_com_tile_module_n_142, ZN => vga_com_tile_module_n_141);
  vga_com_tile_module_g48573 : CKND1BWP7T port map(I => vga_com_tile_module_n_139, ZN => vga_com_tile_module_n_138);
  vga_com_tile_module_g48574 : INVD0BWP7T port map(I => vga_com_tile_module_n_136, ZN => vga_com_tile_module_n_135);
  vga_com_tile_module_g48575 : INVD0BWP7T port map(I => vga_com_tile_module_n_134, ZN => vga_com_tile_module_n_133);
  vga_com_tile_module_g48576 : INVD0BWP7T port map(I => vga_com_tile_module_n_131, ZN => vga_com_tile_module_n_130);
  vga_com_tile_module_g48577 : INVD0BWP7T port map(I => vga_com_tile_module_n_129, ZN => vga_com_tile_module_n_128);
  vga_com_tile_module_g48578 : INVD0BWP7T port map(I => vga_com_tile_module_n_127, ZN => vga_com_tile_module_n_126);
  vga_com_tile_module_g48579 : INVD1BWP7T port map(I => vga_com_tile_module_n_125, ZN => vga_com_tile_module_n_124);
  vga_com_tile_module_g48580 : INVD1BWP7T port map(I => vga_com_tile_module_n_123, ZN => vga_com_tile_module_n_122);
  vga_com_tile_module_g48581 : INVD1BWP7T port map(I => vga_com_tile_module_n_120, ZN => vga_com_tile_module_n_119);
  vga_com_tile_module_g48582 : INVD1BWP7T port map(I => vga_com_tile_module_n_118, ZN => vga_com_tile_module_n_117);
  vga_com_tile_module_g48583 : INVD1BWP7T port map(I => vga_com_tile_module_n_116, ZN => vga_com_tile_module_n_115);
  vga_com_tile_module_g48584 : INVD1BWP7T port map(I => vga_com_tile_module_n_114, ZN => vga_com_tile_module_n_113);
  vga_com_tile_module_g48585 : INVD0BWP7T port map(I => vga_com_tile_module_n_112, ZN => vga_com_tile_module_n_111);
  vga_com_tile_module_g48586 : INVD1BWP7T port map(I => vga_com_tile_module_n_110, ZN => vga_com_tile_module_n_109);
  vga_com_tile_module_g48587 : INVD1BWP7T port map(I => vga_com_tile_module_n_108, ZN => vga_com_tile_module_n_107);
  vga_com_tile_module_g48588 : INVD1BWP7T port map(I => vga_com_tile_module_n_106, ZN => vga_com_tile_module_n_105);
  vga_com_tile_module_g48589 : INVD1BWP7T port map(I => vga_com_tile_module_n_104, ZN => vga_com_tile_module_n_103);
  vga_com_tile_module_g48590 : AOI21D0BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_tile_module_n_4, B => vga_com_tile_module_n_74, ZN => vga_com_tile_module_n_102);
  vga_com_tile_module_g48591 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_85, A2 => vga_com_tile_module_n_65, ZN => vga_com_tile_module_n_176);
  vga_com_tile_module_g48592 : CKND2D0BWP7T port map(A1 => vga_com_tile_module_n_79, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_175);
  vga_com_tile_module_g48593 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_26, A2 => vga_com_tile_module_n_64, ZN => vga_com_tile_module_n_174);
  vga_com_tile_module_g48594 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_66, A2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_173);
  vga_com_tile_module_g48595 : CKXOR2D1BWP7T port map(A1 => vga_com_bg_select(2), A2 => vga_com_bg_select(1), Z => vga_com_tile_module_n_172);
  vga_com_tile_module_g48596 : CKND2D0BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_171);
  vga_com_tile_module_g48597 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_17, A2 => vga_com_tile_module_n_64, ZN => vga_com_tile_module_n_170);
  vga_com_tile_module_g48598 : ND2D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_169);
  vga_com_tile_module_g48599 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_72, A2 => vga_com_tile_module_n_41, ZN => vga_com_tile_module_n_168);
  vga_com_tile_module_g48600 : NR2D0BWP7T port map(A1 => vga_com_tile_module_n_41, A2 => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_167);
  vga_com_tile_module_g48601 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_36, A2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_165);
  vga_com_tile_module_g48602 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_40, A2 => vga_com_tile_module_n_85, ZN => vga_com_tile_module_n_163);
  vga_com_tile_module_g48603 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_2, A2 => vga_com_tile_module_n_57, ZN => vga_com_tile_module_n_162);
  vga_com_tile_module_g48604 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_78, A2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_161);
  vga_com_tile_module_g48605 : NR2D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => vga_com_tile_module_n_53, ZN => vga_com_tile_module_n_160);
  vga_com_tile_module_g48606 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_83, A2 => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_158);
  vga_com_tile_module_g48607 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_2, A2 => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_157);
  vga_com_tile_module_g48608 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_62, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_156);
  vga_com_tile_module_g48609 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_39, A2 => vga_com_tile_module_n_22, ZN => vga_com_tile_module_n_155);
  vga_com_tile_module_g48610 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_36, A2 => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_153);
  vga_com_tile_module_g48611 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_39, A2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_152);
  vga_com_tile_module_g48612 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_33, A2 => vga_com_tile_module_n_22, ZN => vga_com_tile_module_n_150);
  vga_com_tile_module_g48613 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_39, A2 => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_149);
  vga_com_tile_module_g48614 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_39, A2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_147);
  vga_com_tile_module_g48615 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_27, A2 => vga_com_tile_module_n_28, ZN => vga_com_tile_module_n_146);
  vga_com_tile_module_g48616 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_67, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_144);
  vga_com_tile_module_g48617 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_33, A2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_143);
  vga_com_tile_module_g48618 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_35, A2 => vga_com_tile_module_n_21, ZN => vga_com_tile_module_n_142);
  vga_com_tile_module_g48619 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_47, A2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_140);
  vga_com_tile_module_g48620 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_35, A2 => vga_com_tile_module_n_30, ZN => vga_com_tile_module_n_139);
  vga_com_tile_module_g48621 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_35, A2 => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_137);
  vga_com_tile_module_g48622 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_33, A2 => vga_com_tile_module_n_20, ZN => vga_com_tile_module_n_136);
  vga_com_tile_module_g48623 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_36, A2 => vga_com_tile_module_n_20, ZN => vga_com_tile_module_n_134);
  vga_com_tile_module_g48624 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_64, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_132);
  vga_com_tile_module_g48625 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_37, A2 => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_131);
  vga_com_tile_module_g48626 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_34, A2 => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_129);
  vga_com_tile_module_g48627 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_32, A2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_127);
  vga_com_tile_module_g48628 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_33, A2 => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_125);
  vga_com_tile_module_g48629 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_32, A2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_123);
  vga_com_tile_module_g48630 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_51, A2 => vga_com_tile_module_n_64, ZN => vga_com_tile_module_n_121);
  vga_com_tile_module_g48631 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_41, A2 => vga_com_tile_module_n_66, ZN => vga_com_tile_module_n_120);
  vga_com_tile_module_g48632 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_31, A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_118);
  vga_com_tile_module_g48633 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_65, A2 => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_116);
  vga_com_tile_module_g48634 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_31, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_114);
  vga_com_tile_module_g48635 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_25, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_112);
  vga_com_tile_module_g48636 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_17, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_110);
  vga_com_tile_module_g48637 : NR2D1P5BWP7T port map(A1 => vga_com_tile_module_n_35, A2 => vga_com_tile_module_n_10, ZN => vga_com_tile_module_n_108);
  vga_com_tile_module_g48638 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_23, A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_106);
  vga_com_tile_module_g48639 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_25, A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_104);
  vga_com_tile_module_g48640 : INVD1BWP7T port map(I => vga_com_tile_module_n_92, ZN => vga_com_tile_module_n_91);
  vga_com_tile_module_g48641 : INVD0BWP7T port map(I => vga_com_tile_module_n_90, ZN => vga_com_tile_module_n_89);
  vga_com_tile_module_g48642 : INVD0BWP7T port map(I => vga_com_tile_module_n_88, ZN => vga_com_tile_module_n_87);
  vga_com_tile_module_g48643 : INVD0BWP7T port map(I => vga_com_tile_module_n_85, ZN => vga_com_tile_module_n_84);
  vga_com_tile_module_g48644 : INVD1BWP7T port map(I => vga_com_tile_module_n_83, ZN => vga_com_tile_module_n_82);
  vga_com_tile_module_g48645 : INVD1BWP7T port map(I => vga_com_tile_module_n_81, ZN => vga_com_tile_module_n_80);
  vga_com_tile_module_g48646 : INVD1BWP7T port map(I => vga_com_tile_module_n_79, ZN => vga_com_tile_module_n_78);
  vga_com_tile_module_g48647 : INVD1BWP7T port map(I => vga_com_tile_module_n_77, ZN => vga_com_tile_module_n_76);
  vga_com_tile_module_g48648 : INVD1BWP7T port map(I => vga_com_tile_module_n_75, ZN => vga_com_tile_module_n_74);
  vga_com_tile_module_g48649 : INVD1BWP7T port map(I => vga_com_tile_module_n_73, ZN => vga_com_tile_module_n_72);
  vga_com_tile_module_g48650 : INVD1BWP7T port map(I => vga_com_tile_module_n_71, ZN => vga_com_tile_module_n_70);
  vga_com_tile_module_g48651 : INVD1BWP7T port map(I => vga_com_tile_module_n_69, ZN => vga_com_tile_module_n_68);
  vga_com_tile_module_g48652 : INVD1BWP7T port map(I => vga_com_tile_module_n_67, ZN => vga_com_tile_module_n_66);
  vga_com_tile_module_g48653 : INVD1BWP7T port map(I => vga_com_tile_module_n_65, ZN => vga_com_tile_module_n_64);
  vga_com_tile_module_g48654 : INVD1BWP7T port map(I => vga_com_tile_module_n_63, ZN => vga_com_tile_module_n_62);
  vga_com_tile_module_g48655 : CKND2D0BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => vga_com_column(2), ZN => vga_com_tile_module_n_101);
  vga_com_tile_module_g48656 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_7, A2 => vga_com_bg_select(1), ZN => vga_com_tile_module_n_100);
  vga_com_tile_module_g48657 : NR2XD0BWP7T port map(A1 => vga_com_tile_address(5), A2 => FE_OFN0_reset, ZN => vga_com_tile_module_n_99);
  vga_com_tile_module_g48658 : ND2D1BWP7T port map(A1 => vga_com_tile_address(3), A2 => vga_com_tile_address(4), ZN => vga_com_tile_module_n_98);
  vga_com_tile_module_g48659 : ND2D1BWP7T port map(A1 => vga_com_tile_address(3), A2 => vga_com_tile_module_n_13, ZN => vga_com_tile_module_n_97);
  vga_com_tile_module_g48660 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_6, A2 => vga_com_tile_address(4), ZN => vga_com_tile_module_n_96);
  vga_com_tile_module_g48661 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_5, A2 => vga_com_tile_address(3), ZN => vga_com_tile_module_n_95);
  vga_com_tile_module_g48662 : NR2XD0BWP7T port map(A1 => vga_com_tile_address(3), A2 => vga_com_tile_address(4), ZN => vga_com_tile_module_n_94);
  vga_com_tile_module_g48663 : IND2D1BWP7T port map(A1 => FE_OFN0_reset, B1 => vga_com_tile_address(5), ZN => vga_com_tile_module_n_93);
  vga_com_tile_module_g48664 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_92);
  vga_com_tile_module_g48665 : ND2D1BWP7T port map(A1 => vga_com_tile_address(2), A2 => vga_com_tile_address(3), ZN => vga_com_tile_module_n_90);
  vga_com_tile_module_g48666 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_tile_module_n_11, ZN => vga_com_tile_module_n_88);
  vga_com_tile_module_g48667 : NR2D1BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_address(2), ZN => vga_com_tile_module_n_86);
  vga_com_tile_module_g48668 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_column(1), ZN => vga_com_tile_module_n_85);
  vga_com_tile_module_g48669 : ND2D1BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_address(2), ZN => vga_com_tile_module_n_83);
  vga_com_tile_module_g48670 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_tile_module_n_11, ZN => vga_com_tile_module_n_81);
  vga_com_tile_module_g48671 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_column(1), ZN => vga_com_tile_module_n_79);
  vga_com_tile_module_g48672 : CKND2D1BWP7T port map(A1 => vga_com_column(0), A2 => vga_com_column(1), ZN => vga_com_tile_module_n_77);
  vga_com_tile_module_g48673 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_tile_module_n_12, ZN => vga_com_tile_module_n_75);
  vga_com_tile_module_g48674 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_12, A2 => vga_com_column(2), ZN => vga_com_tile_module_n_73);
  vga_com_tile_module_g48675 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_3, A2 => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_71);
  vga_com_tile_module_g48676 : NR2XD0BWP7T port map(A1 => vga_com_tile_address(1), A2 => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_69);
  vga_com_tile_module_g48677 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_11, A2 => vga_com_column(1), ZN => vga_com_tile_module_n_67);
  vga_com_tile_module_g48678 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_11, A2 => vga_com_tile_module_n_12, ZN => vga_com_tile_module_n_65);
  vga_com_tile_module_g48679 : ND2D1BWP7T port map(A1 => vga_com_column(1), A2 => vga_com_column(2), ZN => vga_com_tile_module_n_63);
  vga_com_tile_module_g48680 : INVD1BWP7T port map(I => vga_com_tile_module_n_59, ZN => vga_com_tile_module_n_58);
  vga_com_tile_module_g48681 : INVD0BWP7T port map(I => vga_com_tile_module_n_57, ZN => vga_com_tile_module_n_56);
  vga_com_tile_module_g48682 : INVD1BWP7T port map(I => vga_com_tile_module_n_55, ZN => vga_com_tile_module_n_54);
  vga_com_tile_module_g48683 : INVD1BWP7T port map(I => vga_com_tile_module_n_53, ZN => vga_com_tile_module_n_52);
  vga_com_tile_module_g48684 : INVD1BWP7T port map(I => vga_com_tile_module_n_51, ZN => vga_com_tile_module_n_50);
  vga_com_tile_module_g48685 : CKND1BWP7T port map(I => vga_com_tile_module_n_49, ZN => vga_com_tile_module_n_48);
  vga_com_tile_module_g48686 : INVD0BWP7T port map(I => vga_com_tile_module_n_47, ZN => vga_com_tile_module_n_46);
  vga_com_tile_module_g48687 : INVD1BWP7T port map(I => vga_com_tile_module_n_45, ZN => vga_com_tile_module_n_44);
  vga_com_tile_module_g48688 : INVD1BWP7T port map(I => vga_com_tile_module_n_43, ZN => vga_com_tile_module_n_42);
  vga_com_tile_module_g48689 : INVD1BWP7T port map(I => vga_com_tile_module_n_41, ZN => vga_com_tile_module_n_40);
  vga_com_tile_module_g48690 : INVD1BWP7T port map(I => vga_com_tile_module_n_39, ZN => vga_com_tile_module_n_38);
  vga_com_tile_module_g48691 : INVD1BWP7T port map(I => vga_com_tile_module_n_37, ZN => vga_com_tile_module_n_36);
  vga_com_tile_module_g48692 : INVD1BWP7T port map(I => vga_com_tile_module_n_35, ZN => vga_com_tile_module_n_34);
  vga_com_tile_module_g48693 : INVD1BWP7T port map(I => vga_com_tile_module_n_33, ZN => vga_com_tile_module_n_32);
  vga_com_tile_module_g48694 : INVD1BWP7T port map(I => vga_com_tile_module_n_31, ZN => vga_com_tile_module_n_30);
  vga_com_tile_module_g48695 : INVD1BWP7T port map(I => vga_com_tile_module_n_29, ZN => vga_com_tile_module_n_28);
  vga_com_tile_module_g48696 : INVD1BWP7T port map(I => vga_com_tile_module_n_27, ZN => vga_com_tile_module_n_26);
  vga_com_tile_module_g48697 : INVD1BWP7T port map(I => vga_com_tile_module_n_25, ZN => vga_com_tile_module_n_24);
  vga_com_tile_module_g48698 : INVD1BWP7T port map(I => vga_com_tile_module_n_23, ZN => vga_com_tile_module_n_22);
  vga_com_tile_module_g48699 : INVD1BWP7T port map(I => vga_com_tile_module_n_21, ZN => vga_com_tile_module_n_20);
  vga_com_tile_module_g48700 : INVD1BWP7T port map(I => vga_com_tile_module_n_19, ZN => vga_com_tile_module_n_18);
  vga_com_tile_module_g48701 : INVD1BWP7T port map(I => vga_com_tile_module_n_17, ZN => vga_com_tile_module_n_16);
  vga_com_tile_module_g48702 : ND2D0BWP7T port map(A1 => vga_com_tile_module_n_11, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_15);
  vga_com_tile_module_g48703 : ND2D1BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_61);
  vga_com_tile_module_g48704 : ND2D1BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_60);
  vga_com_tile_module_g48705 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_11, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_59);
  vga_com_tile_module_g48706 : NR2D1BWP7T port map(A1 => FE_OFN1_vga_com_row_0, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_57);
  vga_com_tile_module_g48707 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_3, A2 => vga_com_tile_address(2), ZN => vga_com_tile_module_n_55);
  vga_com_tile_module_g48708 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_9, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_53);
  vga_com_tile_module_g48709 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_51);
  vga_com_tile_module_g48710 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_3, A2 => vga_com_tile_address(2), ZN => vga_com_tile_module_n_49);
  vga_com_tile_module_g48711 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_column(2), ZN => vga_com_tile_module_n_47);
  vga_com_tile_module_g48712 : NR2XD0BWP7T port map(A1 => vga_com_tile_module_n_3, A2 => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_45);
  vga_com_tile_module_g48713 : NR2D1BWP7T port map(A1 => vga_com_tile_address(1), A2 => vga_com_tile_module_n_2, ZN => vga_com_tile_module_n_43);
  vga_com_tile_module_g48714 : NR2D1BWP7T port map(A1 => vga_com_tile_module_n_4, A2 => vga_com_column(2), ZN => vga_com_tile_module_n_41);
  vga_com_tile_module_g48715 : NR2D1P5BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_39);
  vga_com_tile_module_g48716 : ND2D1BWP7T port map(A1 => vga_com_tile_module_n_2, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_37);
  vga_com_tile_module_g48717 : ND2D1BWP7T port map(A1 => FE_OFN2_vga_com_tile_address_0, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_35);
  vga_com_tile_module_g48718 : NR2D1P5BWP7T port map(A1 => vga_com_tile_module_n_2, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_33);
  vga_com_tile_module_g48719 : NR2D1P5BWP7T port map(A1 => vga_com_tile_module_n_8, A2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_31);
  vga_com_tile_module_g48720 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_9, A2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_29);
  vga_com_tile_module_g48721 : NR2D1P5BWP7T port map(A1 => vga_com_tile_module_n_9, A2 => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_27);
  vga_com_tile_module_g48722 : NR2XD1BWP7T port map(A1 => vga_com_tile_module_n_10, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_25);
  vga_com_tile_module_g48723 : CKND2D1BWP7T port map(A1 => FE_OFN3_vga_com_row_1, A2 => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_23);
  vga_com_tile_module_g48724 : CKND2D1BWP7T port map(A1 => vga_com_tile_module_n_10, A2 => vga_com_tile_module_n_8, ZN => vga_com_tile_module_n_21);
  vga_com_tile_module_g48725 : NR2D1P5BWP7T port map(A1 => vga_com_tile_module_n_10, A2 => vga_com_tile_module_n_9, ZN => vga_com_tile_module_n_19);
  vga_com_tile_module_g48726 : NR2D1P5BWP7T port map(A1 => FE_OFN3_vga_com_row_1, A2 => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_17);
  vga_com_tile_module_g48727 : INVD1BWP7T port map(I => vga_com_timer1(5), ZN => vga_com_tile_module_n_14);
  vga_com_tile_module_g48728 : INVD0BWP7T port map(I => vga_com_tile_address(4), ZN => vga_com_tile_module_n_13);
  vga_com_tile_module_g48729 : INVD1BWP7T port map(I => vga_com_column(1), ZN => vga_com_tile_module_n_12);
  vga_com_tile_module_g48730 : INVD1BWP7T port map(I => vga_com_column(2), ZN => vga_com_tile_module_n_11);
  vga_com_tile_module_g48731 : INVD1P5BWP7T port map(I => FE_OFN3_vga_com_row_1, ZN => vga_com_tile_module_n_10);
  vga_com_tile_module_g48732 : INVD1P5BWP7T port map(I => FE_OFN4_vga_com_row_2, ZN => vga_com_tile_module_n_9);
  vga_com_tile_module_g48733 : INVD1BWP7T port map(I => FE_OFN1_vga_com_row_0, ZN => vga_com_tile_module_n_8);
  vga_com_tile_module_g48734 : CKND1BWP7T port map(I => vga_com_bg_select(0), ZN => vga_com_tile_module_n_7);
  vga_com_tile_module_g48735 : INVD1BWP7T port map(I => vga_com_tile_address(3), ZN => vga_com_tile_module_n_6);
  vga_com_tile_module_g48736 : INVD1BWP7T port map(I => vga_com_tile_address(2), ZN => vga_com_tile_module_n_5);
  vga_com_tile_module_g48737 : INVD1BWP7T port map(I => vga_com_column(0), ZN => vga_com_tile_module_n_4);
  vga_com_tile_module_g48738 : INVD1BWP7T port map(I => vga_com_tile_address(1), ZN => vga_com_tile_module_n_3);
  vga_com_tile_module_g48739 : INVD1BWP7T port map(I => FE_OFN2_vga_com_tile_address_0, ZN => vga_com_tile_module_n_2);
  vga_com_tile_module_g2 : OA21D0BWP7T port map(A1 => vga_com_tile_module_n_448, A2 => vga_com_tile_module_n_10, B => vga_com_tile_module_n_462, Z => vga_com_tile_module_n_1);
  vga_com_tile_module_g48740 : IND2D1BWP7T port map(A1 => vga_com_tile_module_n_172, B1 => vga_com_bg_select(0), ZN => vga_com_tile_module_n_0);
  vga_com_tile_module_g48741 : OAI21D0BWP7T port map(A1 => vga_com_tile_module_n_342, A2 => vga_com_tile_module_n_10, B => vga_com_tile_module_n_259, ZN => vga_com_tile_module_n_1060);
  vga_com_color_driver_module_g870 : ND3D0BWP7T port map(A1 => vga_com_color_driver_module_n_55, A2 => vga_com_color_driver_module_n_33, A3 => vga_com_color_driver_module_n_15, ZN => vga_com_in_red(2));
  vga_com_color_driver_module_g871 : ND4D0BWP7T port map(A1 => vga_com_color_driver_module_n_50, A2 => vga_com_color_driver_module_n_40, A3 => vga_com_color_driver_module_n_38, A4 => vga_com_color_driver_module_n_26, ZN => vga_com_in_blue(2));
  vga_com_color_driver_module_g872 : ND4D0BWP7T port map(A1 => vga_com_color_driver_module_n_51, A2 => vga_com_color_driver_module_n_38, A3 => vga_com_color_driver_module_n_37, A4 => vga_com_color_driver_module_n_36, ZN => vga_com_in_blue(3));
  vga_com_color_driver_module_g873 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_52, A2 => vga_com_color_driver_module_n_28, ZN => vga_com_in_red(1));
  vga_com_color_driver_module_g874 : OAI211D1BWP7T port map(A1 => vga_com_color_driver_module_n_6, A2 => vga_com_color_driver_module_n_23, B => vga_com_color_driver_module_n_41, C => vga_com_color_driver_module_n_37, ZN => vga_com_in_green(1));
  vga_com_color_driver_module_g875 : ND3D0BWP7T port map(A1 => vga_com_color_driver_module_n_44, A2 => vga_com_color_driver_module_n_45, A3 => vga_com_color_driver_module_n_26, ZN => vga_com_in_blue(1));
  vga_com_color_driver_module_g876 : AO211D0BWP7T port map(A1 => vga_com_color_driver_module_n_20, A2 => vga_com_color_address(3), B => vga_com_color_driver_module_n_49, C => vga_com_color_driver_module_n_42, Z => vga_com_in_green(2));
  vga_com_color_driver_module_g877 : IND3D1BWP7T port map(A1 => vga_com_color_driver_module_n_43, B1 => vga_com_color_driver_module_n_28, B2 => vga_com_color_driver_module_n_37, ZN => vga_com_in_green(3));
  vga_com_color_driver_module_g878 : AOI222D0BWP7T port map(A1 => vga_com_color_driver_module_n_35, A2 => vga_com_color_address(0), B1 => vga_com_color_driver_module_n_13, B2 => vga_com_color_driver_module_n_8, C1 => vga_com_color_driver_module_n_14, C2 => vga_com_color_address(1), ZN => vga_com_color_driver_module_n_55);
  vga_com_color_driver_module_g879 : AO211D0BWP7T port map(A1 => vga_com_color_driver_module_n_18, A2 => vga_com_color_driver_module_n_13, B => vga_com_color_driver_module_n_49, C => vga_com_color_driver_module_n_31, Z => vga_com_in_red(3));
  vga_com_color_driver_module_g880 : ND3D0BWP7T port map(A1 => vga_com_color_driver_module_n_30, A2 => vga_com_color_driver_module_n_26, A3 => vga_com_color_driver_module_n_19, ZN => vga_com_in_green(0));
  vga_com_color_driver_module_g881 : OA221D0BWP7T port map(A1 => vga_com_color_driver_module_n_25, A2 => vga_com_color_driver_module_n_10, B1 => vga_com_color_address(0), B2 => vga_com_color_driver_module_n_19, C => vga_com_color_driver_module_n_47, Z => vga_com_color_driver_module_n_52);
  vga_com_color_driver_module_g882 : AOI21D0BWP7T port map(A1 => vga_com_color_driver_module_n_34, A2 => vga_com_color_driver_module_n_7, B => vga_com_color_driver_module_n_39, ZN => vga_com_color_driver_module_n_51);
  vga_com_color_driver_module_g883 : AOI32D1BWP7T port map(A1 => vga_com_color_driver_module_n_14, A2 => vga_com_color_driver_module_n_1, A3 => vga_com_color_address(2), B1 => vga_com_color_driver_module_n_34, B2 => vga_com_color_driver_module_n_0, ZN => vga_com_color_driver_module_n_50);
  vga_com_color_driver_module_g884 : ND3D0BWP7T port map(A1 => vga_com_color_driver_module_n_19, A2 => vga_com_color_driver_module_n_29, A3 => vga_com_color_driver_module_n_11, ZN => vga_com_in_red(0));
  vga_com_color_driver_module_g885 : OA21D0BWP7T port map(A1 => vga_com_color_driver_module_n_15, A2 => vga_com_color_driver_module_n_0, B => vga_com_color_driver_module_n_33, Z => vga_com_color_driver_module_n_47);
  vga_com_color_driver_module_g886 : OAI221D0BWP7T port map(A1 => vga_com_color_driver_module_n_7, A2 => vga_com_color_address(4), B1 => vga_com_color_address(2), B2 => vga_com_color_driver_module_n_11, C => vga_com_color_driver_module_n_6, ZN => vga_com_in_blue(0));
  vga_com_color_driver_module_g887 : ND3D0BWP7T port map(A1 => vga_com_color_driver_module_n_21, A2 => vga_com_color_driver_module_n_13, A3 => vga_com_color_address(2), ZN => vga_com_color_driver_module_n_45);
  vga_com_color_driver_module_g888 : OAI21D0BWP7T port map(A1 => vga_com_color_driver_module_n_29, A2 => vga_com_color_address(2), B => vga_com_color_driver_module_n_27, ZN => vga_com_color_driver_module_n_49);
  vga_com_color_driver_module_g889 : OAI21D0BWP7T port map(A1 => vga_com_color_driver_module_n_22, A2 => vga_com_color_driver_module_n_20, B => vga_com_color_driver_module_n_16, ZN => vga_com_color_driver_module_n_44);
  vga_com_color_driver_module_g890 : OAI31D0BWP7T port map(A1 => vga_com_color_address(2), A2 => vga_com_color_driver_module_n_16, A3 => vga_com_color_driver_module_n_12, B => vga_com_color_driver_module_n_32, ZN => vga_com_color_driver_module_n_43);
  vga_com_color_driver_module_g891 : AO22D0BWP7T port map(A1 => vga_com_color_driver_module_n_21, A2 => vga_com_color_driver_module_n_0, B1 => vga_com_color_driver_module_n_1, B2 => vga_com_color_driver_module_n_8, Z => vga_com_color_driver_module_n_42);
  vga_com_color_driver_module_g892 : MAOI22D0BWP7T port map(A1 => vga_com_color_driver_module_n_8, A2 => vga_com_color_address(0), B1 => vga_com_color_driver_module_n_27, B2 => vga_com_color_driver_module_n_12, ZN => vga_com_color_driver_module_n_41);
  vga_com_color_driver_module_g893 : MAOI22D0BWP7T port map(A1 => vga_com_color_driver_module_n_24, A2 => vga_com_color_driver_module_n_10, B1 => vga_com_color_driver_module_n_19, B2 => vga_com_color_driver_module_n_13, ZN => vga_com_color_driver_module_n_40);
  vga_com_color_driver_module_g894 : OAI22D0BWP7T port map(A1 => vga_com_color_driver_module_n_19, A2 => vga_com_color_driver_module_n_7, B1 => vga_com_color_driver_module_n_10, B2 => vga_com_color_driver_module_n_6, ZN => vga_com_color_driver_module_n_39);
  vga_com_color_driver_module_g895 : CKND2D0BWP7T port map(A1 => vga_com_color_driver_module_n_24, A2 => vga_com_color_address(0), ZN => vga_com_color_driver_module_n_36);
  vga_com_color_driver_module_g896 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_28, A2 => vga_com_color_address(3), ZN => vga_com_color_driver_module_n_35);
  vga_com_color_driver_module_g897 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_22, A2 => vga_com_color_driver_module_n_3, ZN => vga_com_color_driver_module_n_38);
  vga_com_color_driver_module_g898 : IND2D1BWP7T port map(A1 => vga_com_color_address(3), B1 => vga_com_color_driver_module_n_20, ZN => vga_com_color_driver_module_n_37);
  vga_com_color_driver_module_g899 : OAI21D0BWP7T port map(A1 => vga_com_color_driver_module_n_4, A2 => vga_com_color_address(1), B => vga_com_color_driver_module_n_21, ZN => vga_com_color_driver_module_n_32);
  vga_com_color_driver_module_g900 : OAI22D0BWP7T port map(A1 => vga_com_color_driver_module_n_0, A2 => vga_com_color_driver_module_n_11, B1 => vga_com_color_driver_module_n_1, B2 => vga_com_color_address(3), ZN => vga_com_color_driver_module_n_31);
  vga_com_color_driver_module_g901 : AOI22D0BWP7T port map(A1 => vga_com_color_driver_module_n_9, A2 => vga_com_color_driver_module_n_8, B1 => vga_com_color_driver_module_n_7, B2 => vga_com_color_driver_module_n_5, ZN => vga_com_color_driver_module_n_30);
  vga_com_color_driver_module_g902 : OAI21D0BWP7T port map(A1 => vga_com_color_driver_module_n_6, A2 => vga_com_color_address(2), B => vga_com_color_driver_module_n_27, ZN => vga_com_color_driver_module_n_34);
  vga_com_color_driver_module_g903 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_20, A2 => vga_com_color_driver_module_n_3, ZN => vga_com_color_driver_module_n_33);
  vga_com_color_driver_module_g904 : CKND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_14, A2 => vga_com_color_address(0), ZN => vga_com_color_driver_module_n_29);
  vga_com_color_driver_module_g905 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_8, A2 => vga_com_color_address(1), ZN => vga_com_color_driver_module_n_28);
  vga_com_color_driver_module_g906 : OR2D1BWP7T port map(A1 => vga_com_color_driver_module_n_15, A2 => vga_com_color_driver_module_n_3, Z => vga_com_color_driver_module_n_27);
  vga_com_color_driver_module_g907 : IND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_7, B1 => vga_com_color_driver_module_n_14, ZN => vga_com_color_driver_module_n_26);
  vga_com_color_driver_module_g908 : INVD1BWP7T port map(I => vga_com_color_driver_module_n_24, ZN => vga_com_color_driver_module_n_25);
  vga_com_color_driver_module_g909 : INVD0BWP7T port map(I => vga_com_color_driver_module_n_22, ZN => vga_com_color_driver_module_n_23);
  vga_com_color_driver_module_g910 : INVD0BWP7T port map(I => vga_com_color_driver_module_n_19, ZN => vga_com_color_driver_module_n_18);
  vga_com_color_driver_module_g911 : NR2XD0BWP7T port map(A1 => vga_com_color_driver_module_n_17, A2 => vga_com_color_address(2), ZN => vga_com_color_driver_module_n_24);
  vga_com_color_driver_module_g912 : NR2XD0BWP7T port map(A1 => vga_com_color_driver_module_n_10, A2 => vga_com_color_address(2), ZN => vga_com_color_driver_module_n_22);
  vga_com_color_driver_module_g913 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_17, A2 => vga_com_color_driver_module_n_6, ZN => vga_com_color_driver_module_n_21);
  vga_com_color_driver_module_g914 : NR2XD0BWP7T port map(A1 => vga_com_color_driver_module_n_7, A2 => vga_com_color_address(2), ZN => vga_com_color_driver_module_n_20);
  vga_com_color_driver_module_g915 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_5, A2 => vga_com_color_address(2), ZN => vga_com_color_driver_module_n_19);
  vga_com_color_driver_module_g916 : INVD0BWP7T port map(I => vga_com_color_driver_module_n_13, ZN => vga_com_color_driver_module_n_12);
  vga_com_color_driver_module_g917 : IND2D1BWP7T port map(A1 => vga_com_color_address(3), B1 => vga_com_color_address(4), ZN => vga_com_color_driver_module_n_17);
  vga_com_color_driver_module_g918 : ND2D1BWP7T port map(A1 => vga_com_color_address(3), A2 => vga_com_color_address(4), ZN => vga_com_color_driver_module_n_16);
  vga_com_color_driver_module_g919 : IND2D1BWP7T port map(A1 => vga_com_color_address(3), B1 => vga_com_color_address(2), ZN => vga_com_color_driver_module_n_15);
  vga_com_color_driver_module_g920 : NR2D1BWP7T port map(A1 => vga_com_color_address(3), A2 => vga_com_color_address(4), ZN => vga_com_color_driver_module_n_14);
  vga_com_color_driver_module_g921 : NR2D1BWP7T port map(A1 => vga_com_color_address(0), A2 => vga_com_color_address(1), ZN => vga_com_color_driver_module_n_13);
  vga_com_color_driver_module_g922 : INVD0BWP7T port map(I => vga_com_color_driver_module_n_10, ZN => vga_com_color_driver_module_n_9);
  vga_com_color_driver_module_g923 : INVD0BWP7T port map(I => vga_com_color_driver_module_n_6, ZN => vga_com_color_driver_module_n_5);
  vga_com_color_driver_module_g924 : NR2D1BWP7T port map(A1 => vga_com_color_address(0), A2 => vga_com_color_driver_module_n_2, ZN => vga_com_color_driver_module_n_4);
  vga_com_color_driver_module_g925 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_3, A2 => vga_com_color_address(1), ZN => vga_com_color_driver_module_n_11);
  vga_com_color_driver_module_g926 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_0, A2 => vga_com_color_address(1), ZN => vga_com_color_driver_module_n_10);
  vga_com_color_driver_module_g927 : NR2D1BWP7T port map(A1 => vga_com_color_driver_module_n_2, A2 => vga_com_color_address(4), ZN => vga_com_color_driver_module_n_8);
  vga_com_color_driver_module_g928 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_1, A2 => vga_com_color_address(0), ZN => vga_com_color_driver_module_n_7);
  vga_com_color_driver_module_g929 : ND2D1BWP7T port map(A1 => vga_com_color_driver_module_n_3, A2 => vga_com_color_address(3), ZN => vga_com_color_driver_module_n_6);
  vga_com_color_driver_module_g930 : INVD1BWP7T port map(I => vga_com_color_address(4), ZN => vga_com_color_driver_module_n_3);
  vga_com_color_driver_module_g931 : INVD0BWP7T port map(I => vga_com_color_address(2), ZN => vga_com_color_driver_module_n_2);
  vga_com_color_driver_module_g932 : INVD1BWP7T port map(I => vga_com_color_address(1), ZN => vga_com_color_driver_module_n_1);
  vga_com_color_driver_module_g933 : INVD1BWP7T port map(I => vga_com_color_address(0), ZN => vga_com_color_driver_module_n_0);
  stable_map_com_map_internal_reg_0 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_90, Q => map_data(0));
  stable_map_com_map_internal_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN258_stable_map_com_n_92, Q => map_data(1));
  stable_map_com_map_internal_reg_2 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_91, Q => map_data(2));
  stable_map_com_map_internal_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_89, Q => map_data(3));
  stable_map_com_map_internal_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_100, Q => map_data(4));
  stable_map_com_map_internal_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN287_stable_map_com_n_111, Q => map_data(5));
  stable_map_com_map_internal_reg_6 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_115, Q => map_data(6));
  stable_map_com_map_internal_reg_7 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_78, Q => map_data(7));
  stable_map_com_map_internal_reg_8 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_85, Q => map_data(8));
  stable_map_com_map_internal_reg_9 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_81, Q => map_data(9));
  stable_map_com_map_internal_reg_10 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_77, Q => map_data(10));
  stable_map_com_map_internal_reg_11 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_74, Q => map_data(11));
  stable_map_com_map_internal_reg_12 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN274_stable_map_com_n_73, Q => map_data(12));
  stable_map_com_map_internal_reg_13 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN293_stable_map_com_n_72, Q => map_data(13));
  stable_map_com_map_internal_reg_14 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN276_stable_map_com_n_71, Q => map_data(14));
  stable_map_com_map_internal_reg_15 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_70, Q => map_data(15));
  stable_map_com_map_internal_reg_16 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_69, Q => map_data(16));
  stable_map_com_map_internal_reg_17 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_67, Q => map_data(17));
  stable_map_com_map_internal_reg_19 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_129, Q => map_data(19));
  stable_map_com_map_internal_reg_20 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_128, Q => map_data(20));
  stable_map_com_map_internal_reg_21 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_105, Q => map_data(21));
  stable_map_com_map_internal_reg_22 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_103, Q => map_data(22));
  stable_map_com_map_internal_reg_23 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_102, Q => map_data(23));
  stable_map_com_map_internal_reg_24 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_101, Q => map_data(24));
  stable_map_com_map_internal_reg_25 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_116, Q => map_data(25));
  stable_map_com_map_internal_reg_26 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_99, Q => map_data(26));
  stable_map_com_map_internal_reg_27 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN289_stable_map_com_n_98, Q => map_data(27));
  stable_map_com_map_internal_reg_28 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_97, Q => map_data(28));
  stable_map_com_map_internal_reg_29 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_96, Q => map_data(29));
  stable_map_com_map_internal_reg_30 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_95, Q => FE_PHN506_map_data_30);
  stable_map_com_map_internal_reg_31 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_94, Q => map_data(31));
  stable_map_com_map_internal_reg_32 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_93, Q => map_data(32));
  stable_map_com_map_internal_reg_33 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN328_stable_map_com_n_136, Q => map_data(33));
  stable_map_com_map_internal_reg_34 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN310_stable_map_com_n_126, Q => map_data(34));
  stable_map_com_map_internal_reg_35 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN278_stable_map_com_n_135, Q => map_data(35));
  stable_map_com_map_internal_reg_37 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN349_stable_map_com_n_130, Q => map_data(37));
  stable_map_com_map_internal_reg_38 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN271_stable_map_com_n_127, Q => map_data(38));
  stable_map_com_map_internal_reg_39 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_112, Q => map_data(39));
  stable_map_com_map_internal_reg_40 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_113, Q => map_data(40));
  stable_map_com_map_internal_reg_41 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_88, Q => map_data(41));
  stable_map_com_map_internal_reg_42 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_87, Q => map_data(42));
  stable_map_com_map_internal_reg_43 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN508_stable_map_com_n_86, Q => map_data(43));
  stable_map_com_map_internal_reg_44 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN471_stable_map_com_n_84, Q => map_data(44));
  stable_map_com_map_internal_reg_45 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_83, Q => map_data(45));
  stable_map_com_map_internal_reg_46 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_82, Q => map_data(46));
  stable_map_com_map_internal_reg_47 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_80, Q => map_data(47));
  stable_map_com_map_internal_reg_48 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN492_stable_map_com_n_79, Q => map_data(48));
  stable_map_com_map_internal_reg_49 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN285_stable_map_com_n_76, Q => map_data(49));
  stable_map_com_map_internal_reg_50 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_75, Q => map_data(50));
  stable_map_com_map_internal_reg_51 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_138, Q => map_data(51));
  stable_map_com_map_internal_reg_52 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN305_stable_map_com_n_137, Q => map_data(52));
  stable_map_com_map_internal_reg_54 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_68, Q => map_data(54));
  stable_map_com_map_internal_reg_55 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_66, Q => map_data(55));
  stable_map_com_map_internal_reg_56 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_65, Q => FE_PHN509_map_data_56);
  stable_map_com_map_internal_reg_57 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_64, Q => map_data(57));
  stable_map_com_map_internal_reg_58 : DFQD1BWP7T port map(CP => CTS_21, D => stable_map_com_n_63, Q => map_data(58));
  stable_map_com_map_internal_reg_59 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_62, Q => map_data(59));
  stable_map_com_map_internal_reg_60 : DFQD1BWP7T port map(CP => CTS_22, D => stable_map_com_n_61, Q => map_data(60));
  stable_map_com_map_internal_reg_61 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN307_stable_map_com_n_60, Q => map_data(61));
  stable_map_com_map_internal_reg_62 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN347_stable_map_com_n_59, Q => map_data(62));
  stable_map_com_map_internal_reg_63 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN427_stable_map_com_n_58, Q => map_data(63));
  stable_map_com_map_internal_reg_64 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_57, Q => FE_PHN457_map_data_64);
  stable_map_com_map_internal_reg_65 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN272_stable_map_com_n_56, Q => map_data(65));
  stable_map_com_map_internal_reg_66 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN332_stable_map_com_n_55, Q => map_data(66));
  stable_map_com_map_internal_reg_67 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN297_stable_map_com_n_109, Q => map_data(67));
  stable_map_com_map_internal_reg_68 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN280_stable_map_com_n_108, Q => map_data(68));
  stable_map_com_map_internal_reg_69 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN346_stable_map_com_n_107, Q => map_data(69));
  stable_map_com_map_internal_reg_70 : DFQD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_106, Q => map_data(70));
  stable_map_com_map_internal_reg_71 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN257_stable_map_com_n_104, Q => map_data(71));
  stable_map_com_state_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => stable_map_com_n_49, Q => stable_map_com_state(0));
  stable_map_com_state_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => stable_map_com_n_121, Q => stable_map_com_state(1));
  stable_map_com_g5434 : ND2D1BWP7T port map(A1 => stable_map_com_n_131, A2 => stable_map_com_n_42, ZN => FE_PHN267_stable_map_com_n_139);
  stable_map_com_g5435 : ND2D1BWP7T port map(A1 => stable_map_com_n_132, A2 => stable_map_com_n_42, ZN => FE_PHN263_stable_map_com_n_138);
  stable_map_com_g5436 : AO222D0BWP7T port map(A1 => stable_map_com_n_125, A2 => map_data(52), B1 => stable_map_com_n_114, B2 => map_data(19), C1 => stable_map_com_n_31, C2 => map_data_volatile(52), Z => stable_map_com_n_137);
  stable_map_com_g5443 : AO221D0BWP7T port map(A1 => stable_map_com_n_117, A2 => map_data(33), B1 => stable_map_com_n_31, B2 => map_data_volatile(33), C => stable_map_com_n_44, Z => stable_map_com_n_136);
  stable_map_com_g5444 : AO221D0BWP7T port map(A1 => stable_map_com_n_117, A2 => map_data(35), B1 => stable_map_com_n_31, B2 => map_data_volatile(35), C => stable_map_com_n_44, Z => stable_map_com_n_135);
  stable_map_com_g5445 : AO22D0BWP7T port map(A1 => stable_map_com_n_122, A2 => map_data(36), B1 => map_data_volatile(36), B2 => stable_map_com_n_31, Z => stable_map_com_n_134);
  stable_map_com_g5446 : AO22D0BWP7T port map(A1 => stable_map_com_n_123, A2 => map_data(18), B1 => map_data_volatile(18), B2 => stable_map_com_n_31, Z => stable_map_com_n_133);
  stable_map_com_g5447 : AOI222D0BWP7T port map(A1 => stable_map_com_n_125, A2 => map_data(51), B1 => stable_map_com_n_52, B2 => map_data(18), C1 => stable_map_com_n_31, C2 => map_data_volatile(51), ZN => stable_map_com_n_132);
  stable_map_com_g5448 : AOI222D0BWP7T port map(A1 => stable_map_com_n_125, A2 => map_data(53), B1 => stable_map_com_n_52, B2 => map_data(20), C1 => stable_map_com_n_31, C2 => map_data_volatile(53), ZN => stable_map_com_n_131);
  stable_map_com_g5449 : IOA21D1BWP7T port map(A1 => stable_map_com_n_31, A2 => FE_PHN181_map_data_volatile_37, B => stable_map_com_n_120, ZN => stable_map_com_n_130);
  stable_map_com_g5450 : IOA21D1BWP7T port map(A1 => stable_map_com_n_31, A2 => FE_PHN43_map_data_volatile_19, B => stable_map_com_n_124, ZN => FE_PHN283_stable_map_com_n_129);
  stable_map_com_g5452 : AO222D0BWP7T port map(A1 => stable_map_com_n_118, A2 => map_data(20), B1 => stable_map_com_n_31, B2 => map_data_volatile(20), C1 => stable_map_com_n_33, C2 => map_data(18), Z => FE_PHN268_stable_map_com_n_128);
  stable_map_com_g5453 : AO222D0BWP7T port map(A1 => stable_map_com_n_119, A2 => map_data(38), B1 => stable_map_com_n_31, B2 => map_data_volatile(38), C1 => stable_map_com_n_36, C2 => map_data(36), Z => stable_map_com_n_127);
  stable_map_com_g5454 : AO22D0BWP7T port map(A1 => stable_map_com_n_110, A2 => map_data(34), B1 => map_data_volatile(34), B2 => stable_map_com_n_31, Z => stable_map_com_n_126);
  stable_map_com_g5488 : OAI21D0BWP7T port map(A1 => stable_map_com_n_53, A2 => stable_map_com_n_46, B => map_data(19), ZN => stable_map_com_n_124);
  stable_map_com_g5489 : OR2D1BWP7T port map(A1 => stable_map_com_n_118, A2 => stable_map_com_n_33, Z => stable_map_com_n_123);
  stable_map_com_g5490 : OR2D1BWP7T port map(A1 => stable_map_com_n_119, A2 => stable_map_com_n_36, Z => stable_map_com_n_122);
  stable_map_com_g5491 : OAI211D1BWP7T port map(A1 => stable_map_com_n_19, A2 => stable_map_com_n_45, B => stable_map_com_n_30, C => FE_DBTN0_reset, ZN => stable_map_com_n_121);
  stable_map_com_g5492 : OAI21D0BWP7T port map(A1 => stable_map_com_n_54, A2 => stable_map_com_n_47, B => map_data(37), ZN => stable_map_com_n_120);
  stable_map_com_g5520 : ND3D0BWP7T port map(A1 => stable_map_com_n_48, A2 => stable_map_com_n_22, A3 => stable_map_com_n_24, ZN => stable_map_com_n_125);
  stable_map_com_g5521 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN493_map_data_25, B1 => map_data_volatile(25), B2 => stable_map_com_n_31, Z => stable_map_com_n_116);
  stable_map_com_g5522 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN411_map_data_6, B1 => FE_PHN94_map_data_volatile_6, B2 => stable_map_com_n_31, Z => stable_map_com_n_115);
  stable_map_com_g5523 : AOI21D0BWP7T port map(A1 => stable_map_com_n_39, A2 => stable_map_com_n_20, B => stable_map_com_n_41, ZN => stable_map_com_n_114);
  stable_map_com_g5524 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN466_map_data_40, B1 => map_data_volatile(40), B2 => stable_map_com_n_31, Z => stable_map_com_n_113);
  stable_map_com_g5525 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN473_map_data_39, B1 => map_data_volatile(39), B2 => stable_map_com_n_31, Z => stable_map_com_n_112);
  stable_map_com_g5526 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(5), B1 => map_data_volatile(5), B2 => stable_map_com_n_31, Z => stable_map_com_n_111);
  stable_map_com_g5527 : OAI21D0BWP7T port map(A1 => stable_map_com_n_38, A2 => stable_map_com_n_16, B => stable_map_com_n_50, ZN => stable_map_com_n_110);
  stable_map_com_g5528 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(67), B1 => FE_PHN60_map_data_volatile_67, B2 => stable_map_com_n_31, Z => stable_map_com_n_109);
  stable_map_com_g5529 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(68), B1 => map_data_volatile(68), B2 => stable_map_com_n_31, Z => stable_map_com_n_108);
  stable_map_com_g5530 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(69), B1 => map_data_volatile(69), B2 => stable_map_com_n_31, Z => stable_map_com_n_107);
  stable_map_com_g5531 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(70), B1 => map_data_volatile(70), B2 => stable_map_com_n_31, Z => FE_PHN350_stable_map_com_n_106);
  stable_map_com_g5532 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN476_map_data_21, B1 => map_data_volatile(21), B2 => stable_map_com_n_31, Z => stable_map_com_n_105);
  stable_map_com_g5533 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(71), B1 => map_data_volatile(71), B2 => stable_map_com_n_31, Z => stable_map_com_n_104);
  stable_map_com_g5534 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN467_map_data_22, B1 => map_data_volatile(22), B2 => stable_map_com_n_31, Z => stable_map_com_n_103);
  stable_map_com_g5535 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(23), B1 => map_data_volatile(23), B2 => stable_map_com_n_31, Z => FE_PHN460_stable_map_com_n_102);
  stable_map_com_g5536 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN464_map_data_24, B1 => FE_PHN74_map_data_volatile_24, B2 => stable_map_com_n_31, Z => stable_map_com_n_101);
  stable_map_com_g5537 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN414_map_data_4, B1 => map_data_volatile(4), B2 => stable_map_com_n_31, Z => stable_map_com_n_100);
  stable_map_com_g5538 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN423_map_data_26, B1 => FE_PHN63_map_data_volatile_26, B2 => stable_map_com_n_31, Z => stable_map_com_n_99);
  stable_map_com_g5539 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(27), B1 => FE_PHN41_map_data_volatile_27, B2 => stable_map_com_n_31, Z => stable_map_com_n_98);
  stable_map_com_g5540 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN486_map_data_28, B1 => FE_PHN47_map_data_volatile_28, B2 => stable_map_com_n_31, Z => stable_map_com_n_97);
  stable_map_com_g5541 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN491_map_data_29, B1 => map_data_volatile(29), B2 => stable_map_com_n_31, Z => stable_map_com_n_96);
  stable_map_com_g5542 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN482_map_data_30, B1 => map_data_volatile(30), B2 => stable_map_com_n_31, Z => stable_map_com_n_95);
  stable_map_com_g5543 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN440_map_data_31, B1 => map_data_volatile(31), B2 => stable_map_com_n_31, Z => stable_map_com_n_94);
  stable_map_com_g5544 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN499_map_data_32, B1 => map_data_volatile(32), B2 => stable_map_com_n_31, Z => stable_map_com_n_93);
  stable_map_com_g5545 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(1), B1 => map_data_volatile(1), B2 => stable_map_com_n_31, Z => stable_map_com_n_92);
  stable_map_com_g5546 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN415_map_data_2, B1 => map_data_volatile(2), B2 => stable_map_com_n_31, Z => stable_map_com_n_91);
  stable_map_com_g5547 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(0), B1 => FE_PHN95_map_data_volatile_0, B2 => stable_map_com_n_31, Z => FE_PHN284_stable_map_com_n_90);
  stable_map_com_g5548 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN438_map_data_3, B1 => map_data_volatile(3), B2 => stable_map_com_n_31, Z => stable_map_com_n_89);
  stable_map_com_g5549 : AO21D0BWP7T port map(A1 => stable_map_com_n_21, A2 => map_data(37), B => stable_map_com_n_54, Z => stable_map_com_n_119);
  stable_map_com_g5550 : AO21D0BWP7T port map(A1 => stable_map_com_n_23, A2 => map_data(19), B => stable_map_com_n_53, Z => stable_map_com_n_118);
  stable_map_com_g5551 : IOA21D1BWP7T port map(A1 => stable_map_com_n_26, A2 => map_data(34), B => stable_map_com_n_50, ZN => stable_map_com_n_117);
  stable_map_com_g5554 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN470_map_data_41, B1 => FE_PHN122_map_data_volatile_41, B2 => stable_map_com_n_31, Z => stable_map_com_n_88);
  stable_map_com_g5555 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN426_map_data_42, B1 => map_data_volatile(42), B2 => stable_map_com_n_31, Z => stable_map_com_n_87);
  stable_map_com_g5556 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN468_map_data_43, B1 => map_data_volatile(43), B2 => stable_map_com_n_31, Z => stable_map_com_n_86);
  stable_map_com_g5557 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN461_map_data_8, B1 => map_data_volatile(8), B2 => stable_map_com_n_31, Z => stable_map_com_n_85);
  stable_map_com_g5558 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(44), B1 => map_data_volatile(44), B2 => stable_map_com_n_31, Z => FE_PHN393_stable_map_com_n_84);
  stable_map_com_g5559 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN469_map_data_45, B1 => map_data_volatile(45), B2 => stable_map_com_n_31, Z => stable_map_com_n_83);
  stable_map_com_g5560 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(46), B1 => FE_PHN179_map_data_volatile_46, B2 => stable_map_com_n_31, Z => FE_PHN345_stable_map_com_n_82);
  stable_map_com_g5561 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN510_map_data_9, B1 => map_data_volatile(9), B2 => stable_map_com_n_31, Z => stable_map_com_n_81);
  stable_map_com_g5562 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN484_map_data_47, B1 => map_data_volatile(47), B2 => stable_map_com_n_31, Z => stable_map_com_n_80);
  stable_map_com_g5563 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(48), B1 => map_data_volatile(48), B2 => stable_map_com_n_31, Z => stable_map_com_n_79);
  stable_map_com_g5564 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(7), B1 => FE_PHN52_map_data_volatile_7, B2 => stable_map_com_n_31, Z => FE_PHN273_stable_map_com_n_78);
  stable_map_com_g5565 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN171_map_data_10, B1 => map_data_volatile(10), B2 => stable_map_com_n_31, Z => stable_map_com_n_77);
  stable_map_com_g5566 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(49), B1 => map_data_volatile(49), B2 => stable_map_com_n_31, Z => stable_map_com_n_76);
  stable_map_com_g5567 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN478_map_data_50, B1 => map_data_volatile(50), B2 => stable_map_com_n_31, Z => stable_map_com_n_75);
  stable_map_com_g5568 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN439_map_data_11, B1 => map_data_volatile(11), B2 => stable_map_com_n_31, Z => stable_map_com_n_74);
  stable_map_com_g5569 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(12), B1 => map_data_volatile(12), B2 => stable_map_com_n_31, Z => stable_map_com_n_73);
  stable_map_com_g5570 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(13), B1 => map_data_volatile(13), B2 => stable_map_com_n_31, Z => stable_map_com_n_72);
  stable_map_com_g5571 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(14), B1 => map_data_volatile(14), B2 => stable_map_com_n_31, Z => stable_map_com_n_71);
  stable_map_com_g5572 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN496_map_data_15, B1 => map_data_volatile(15), B2 => stable_map_com_n_31, Z => stable_map_com_n_70);
  stable_map_com_g5573 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN500_map_data_16, B1 => map_data_volatile(16), B2 => stable_map_com_n_31, Z => stable_map_com_n_69);
  stable_map_com_g5574 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(54), B1 => FE_PHN84_map_data_volatile_54, B2 => stable_map_com_n_31, Z => FE_PHN270_stable_map_com_n_68);
  stable_map_com_g5575 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(17), B1 => FE_PHN61_map_data_volatile_17, B2 => stable_map_com_n_31, Z => FE_PHN277_stable_map_com_n_67);
  stable_map_com_g5576 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN485_map_data_55, B1 => map_data_volatile(55), B2 => stable_map_com_n_31, Z => stable_map_com_n_66);
  stable_map_com_g5577 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN480_map_data_56, B1 => FE_PHN126_map_data_volatile_56, B2 => stable_map_com_n_31, Z => stable_map_com_n_65);
  stable_map_com_g5578 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(57), B1 => map_data_volatile(57), B2 => stable_map_com_n_31, Z => stable_map_com_n_64);
  stable_map_com_g5579 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN416_map_data_58, B1 => map_data_volatile(58), B2 => stable_map_com_n_31, Z => stable_map_com_n_63);
  stable_map_com_g5580 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN483_map_data_59, B1 => FE_PHN45_map_data_volatile_59, B2 => stable_map_com_n_31, Z => stable_map_com_n_62);
  stable_map_com_g5581 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN472_map_data_60, B1 => map_data_volatile(60), B2 => stable_map_com_n_31, Z => stable_map_com_n_61);
  stable_map_com_g5582 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(61), B1 => map_data_volatile(61), B2 => stable_map_com_n_31, Z => stable_map_com_n_60);
  stable_map_com_g5583 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN387_map_data_62, B1 => map_data_volatile(62), B2 => stable_map_com_n_31, Z => stable_map_com_n_59);
  stable_map_com_g5584 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(63), B1 => map_data_volatile(63), B2 => stable_map_com_n_31, Z => stable_map_com_n_58);
  stable_map_com_g5585 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => FE_PHN394_map_data_64, B1 => FE_PHN39_map_data_volatile_64, B2 => stable_map_com_n_31, Z => stable_map_com_n_57);
  stable_map_com_g5586 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(65), B1 => FE_PHN33_map_data_volatile_65, B2 => stable_map_com_n_31, Z => stable_map_com_n_56);
  stable_map_com_g5587 : AO22D0BWP7T port map(A1 => stable_map_com_n_40, A2 => map_data(66), B1 => FE_PHN70_map_data_volatile_66, B2 => stable_map_com_n_31, Z => stable_map_com_n_55);
  stable_map_com_g5588 : NR2XD0BWP7T port map(A1 => stable_map_com_n_45, A2 => stable_map_com_n_10, ZN => stable_map_com_n_51);
  stable_map_com_g5589 : OAI211D1BWP7T port map(A1 => stable_map_com_n_22, A2 => vga_done, B => stable_map_com_n_219, C => stable_map_com_n_24, ZN => stable_map_com_n_54);
  stable_map_com_g5590 : OAI211D1BWP7T port map(A1 => stable_map_com_n_24, A2 => vga_done, B => stable_map_com_n_219, C => stable_map_com_n_22, ZN => stable_map_com_n_53);
  stable_map_com_g5591 : AOI21D0BWP7T port map(A1 => stable_map_com_n_20, A2 => stable_map_com_n_29, B => stable_map_com_n_41, ZN => stable_map_com_n_52);
  stable_map_com_g5592 : OAI22D0BWP7T port map(A1 => stable_map_com_n_28, A2 => vga_done, B1 => stable_map_com_n_18, B2 => stable_map_com_n_34, ZN => FE_PHN338_stable_map_com_n_49);
  stable_map_com_g5593 : INR3D0BWP7T port map(A1 => stable_map_com_n_38, B1 => stable_map_com_n_27, B2 => stable_map_com_n_35, ZN => stable_map_com_n_48);
  stable_map_com_g5594 : OAI31D0BWP7T port map(A1 => map_data(38), A2 => stable_map_com_n_4, A3 => stable_map_com_n_22, B => stable_map_com_n_43, ZN => stable_map_com_n_47);
  stable_map_com_g5595 : OAI32D1BWP7T port map(A1 => map_data(20), A2 => stable_map_com_n_2, A3 => stable_map_com_n_24, B1 => map_data(18), B2 => stable_map_com_n_32, ZN => stable_map_com_n_46);
  stable_map_com_g5596 : NR4D0BWP7T port map(A1 => stable_map_com_n_27, A2 => stable_map_com_n_25, A3 => stable_map_com_n_21, A4 => stable_map_com_n_23, ZN => stable_map_com_n_50);
  stable_map_com_g5597 : ND2D1BWP7T port map(A1 => stable_map_com_n_36, A2 => stable_map_com_n_4, ZN => stable_map_com_n_43);
  stable_map_com_g5598 : IND3D1BWP7T port map(A1 => map_updated, B1 => FE_PHN176_stable_map_com_n_35, B2 => dir_mined(2), ZN => stable_map_com_n_45);
  stable_map_com_g5599 : AN3D0BWP7T port map(A1 => stable_map_com_n_26, A2 => map_data(33), A3 => map_data(35), Z => stable_map_com_n_44);
  stable_map_com_g5600 : AOI31D0BWP7T port map(A1 => stable_map_com_n_9, A2 => stable_map_com_n_12, A3 => map_data(53), B => stable_map_com_n_17, ZN => stable_map_com_n_39);
  stable_map_com_g5601 : IND3D1BWP7T port map(A1 => stable_map_com_n_12, B1 => map_data(53), B2 => stable_map_com_n_25, ZN => stable_map_com_n_42);
  stable_map_com_g5602 : ND3D0BWP7T port map(A1 => vga_done, A2 => stable_map_com_n_25, A3 => stable_map_com_state(2), ZN => stable_map_com_n_41);
  stable_map_com_g5603 : OA31D2BWP7T port map(A1 => stable_map_com_n_11, A2 => stable_map_com_n_13, A3 => stable_map_com_n_8, B => stable_map_com_n_30, Z => stable_map_com_n_40);
  stable_map_com_g5604 : INVD0BWP7T port map(I => FE_PHN176_stable_map_com_n_35, ZN => stable_map_com_n_34);
  stable_map_com_g5605 : ND2D1BWP7T port map(A1 => stable_map_com_n_26, A2 => stable_map_com_state(0), ZN => stable_map_com_n_38);
  stable_map_com_g5607 : INR2D1BWP7T port map(A1 => map_data(38), B1 => stable_map_com_n_22, ZN => stable_map_com_n_36);
  stable_map_com_g5608 : INR2D1BWP7T port map(A1 => stable_map_com_n_25, B1 => stable_map_com_state(2), ZN => stable_map_com_n_35);
  stable_map_com_g5609 : INVD1BWP7T port map(I => stable_map_com_n_32, ZN => stable_map_com_n_33);
  stable_map_com_g5610 : INVD0BWP7T port map(I => stable_map_com_n_31, ZN => stable_map_com_n_30);
  stable_map_com_g5611 : IOA21D0BWP7T port map(A1 => stable_map_com_n_12, A2 => stable_map_com_n_1, B => stable_map_com_n_9, ZN => stable_map_com_n_29);
  stable_map_com_g5612 : AOI22D0BWP7T port map(A1 => stable_map_com_n_8, A2 => stable_map_com_n_7, B1 => stable_map_com_n_13, B2 => stable_map_com_n_3, ZN => stable_map_com_n_28);
  stable_map_com_g5613 : ND2D1BWP7T port map(A1 => stable_map_com_n_23, A2 => map_data(20), ZN => stable_map_com_n_32);
  stable_map_com_g5614 : AN3D2BWP7T port map(A1 => vga_done, A2 => stable_map_com_n_14, A3 => stable_map_com_n_11, Z => stable_map_com_n_31);
  stable_map_com_g5615 : INVD1BWP7T port map(I => stable_map_com_n_24, ZN => stable_map_com_n_23);
  stable_map_com_g5616 : INVD0BWP7T port map(I => stable_map_com_n_22, ZN => stable_map_com_n_21);
  stable_map_com_g5617 : INR2D1BWP7T port map(A1 => stable_map_com_n_11, B1 => vga_done, ZN => stable_map_com_n_27);
  stable_map_com_g5618 : AN2D1BWP7T port map(A1 => stable_map_com_n_11, A2 => stable_map_com_state(2), Z => stable_map_com_n_26);
  stable_map_com_g5619 : INR2D1BWP7T port map(A1 => stable_map_com_n_11, B1 => stable_map_com_state(0), ZN => stable_map_com_n_25);
  stable_map_com_g5620 : ND2D1BWP7T port map(A1 => stable_map_com_n_13, A2 => stable_map_com_state(1), ZN => stable_map_com_n_24);
  stable_map_com_g5621 : ND2D1BWP7T port map(A1 => stable_map_com_n_8, A2 => stable_map_com_state(1), ZN => stable_map_com_n_22);
  stable_map_com_g5622 : AOI21D0BWP7T port map(A1 => dir_mined(1), A2 => dir_mined(0), B => stable_map_com_n_10, ZN => stable_map_com_n_19);
  stable_map_com_g5623 : AOI21D0BWP7T port map(A1 => dir_mined(2), A2 => stable_map_com_n_6, B => map_updated, ZN => stable_map_com_n_18);
  stable_map_com_g5624 : NR2D0BWP7T port map(A1 => stable_map_com_n_12, A2 => map_data(53), ZN => stable_map_com_n_17);
  stable_map_com_g5625 : XNR2D1BWP7T port map(A1 => map_data(33), A2 => map_data(35), ZN => stable_map_com_n_16);
  stable_map_com_g5626 : OR2D1BWP7T port map(A1 => stable_map_com_n_9, A2 => map_data(53), Z => stable_map_com_n_20);
  stable_map_com_g5628 : INR2XD0BWP7T port map(A1 => stable_map_com_state(0), B1 => stable_map_com_state(2), ZN => stable_map_com_n_14);
  stable_map_com_g5629 : AN2D1BWP7T port map(A1 => stable_map_com_state(0), A2 => FE_DBTN0_reset, Z => stable_map_com_n_13);
  stable_map_com_g5630 : CKND2D1BWP7T port map(A1 => map_data(51), A2 => map_data(52), ZN => stable_map_com_n_12);
  stable_map_com_g5631 : NR2XD0BWP7T port map(A1 => stable_map_com_state(1), A2 => FE_OFN0_reset, ZN => stable_map_com_n_11);
  stable_map_com_g5632 : ND2D1BWP7T port map(A1 => stable_map_com_state(0), A2 => stable_map_com_state(1), ZN => stable_map_com_n_7);
  stable_map_com_g5633 : NR2D1BWP7T port map(A1 => dir_mined(1), A2 => dir_mined(0), ZN => stable_map_com_n_10);
  stable_map_com_g5634 : OR2D1BWP7T port map(A1 => map_data(52), A2 => map_data(51), Z => stable_map_com_n_9);
  stable_map_com_g5635 : NR2XD0BWP7T port map(A1 => stable_map_com_n_3, A2 => FE_OFN0_reset, ZN => stable_map_com_n_8);
  stable_map_com_g5636 : INVD0BWP7T port map(I => dir_mined(0), ZN => stable_map_com_n_6);
  stable_map_com_map_internal_reg_36 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN348_stable_map_com_n_134, Q => map_data(36), QN => stable_map_com_n_4);
  stable_map_com_state_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => stable_map_com_n_51, Q => stable_map_com_state(2), QN => stable_map_com_n_3);
  stable_map_com_map_internal_reg_18 : DFD1BWP7T port map(CP => CTS_21, D => FE_PHN323_stable_map_com_n_133, Q => map_data(18), QN => stable_map_com_n_2);
  stable_map_com_map_internal_reg_53 : DFD1BWP7T port map(CP => CTS_20, D => stable_map_com_n_139, Q => map_data(53), QN => stable_map_com_n_1);
  stable_map_com_g2 : IOA21D1BWP7T port map(A1 => vga_done, A2 => stable_map_com_n_14, B => stable_map_com_n_11, ZN => stable_map_com_n_219);
  spi_com_send_in1_reg : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN66_spi_com_send_in0, Q => spi_com_send_in1);
  spi_com_g5923 : CKAN2D8BWP7T port map(A1 => spi_com_n_3, A2 => spi_com_state(1), Z => SCLK);
  spi_com_g5924 : CKAN2D8BWP7T port map(A1 => spi_com_n_3, A2 => spi_com_n_264, Z => SS);
  spi_com_MISO_shift_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN255_spi_com_n_262, Q => FE_PHN144_spi_com_MISO_shift_0);
  spi_com_MISO_shift_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_211, Q => FE_PHN135_spi_com_MISO_shift_1);
  spi_com_MISO_shift_reg_2 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_206, Q => FE_PHN18_spi_com_MISO_shift_2);
  spi_com_MISO_shift_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_203, Q => FE_PHN162_spi_com_MISO_shift_3);
  spi_com_MISO_shift_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_201, Q => FE_PHN46_spi_com_MISO_shift_4);
  spi_com_MISO_shift_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_198, Q => spi_com_MISO_shift(5));
  spi_com_MISO_shift_reg_6 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_235, Q => FE_PHN64_spi_com_MISO_shift_6);
  spi_com_MISO_shift_reg_7 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_172, Q => FE_PHN22_spi_com_MISO_shift_7);
  spi_com_MISO_shift_reg_8 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_192, Q => spi_com_MISO_shift(8));
  spi_com_MISO_shift_reg_9 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_189, Q => FE_PHN97_spi_com_MISO_shift_9);
  spi_com_MISO_shift_reg_10 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_184, Q => FE_PHN68_spi_com_MISO_shift_10);
  spi_com_MISO_shift_reg_11 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN261_spi_com_n_182, Q => FE_PHN173_spi_com_MISO_shift_11);
  spi_com_MISO_shift_reg_12 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_178, Q => spi_com_MISO_shift(12));
  spi_com_MISO_shift_reg_13 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN265_spi_com_n_175, Q => FE_PHN140_spi_com_MISO_shift_13);
  spi_com_MISO_shift_reg_14 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_171, Q => spi_com_MISO_shift(14));
  spi_com_MISO_shift_reg_15 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_170, Q => spi_com_MISO_shift(15));
  spi_com_MISO_shift_reg_16 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_166, Q => spi_com_MISO_shift(16));
  spi_com_MISO_shift_reg_17 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_164, Q => FE_PHN121_spi_com_MISO_shift_17);
  spi_com_MISO_shift_reg_18 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_160, Q => FE_PHN421_spi_com_MISO_shift_18);
  spi_com_MISO_shift_reg_19 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_156, Q => FE_PHN34_spi_com_MISO_shift_19);
  spi_com_MISO_shift_reg_20 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_154, Q => FE_PHN72_spi_com_MISO_shift_20);
  spi_com_MISO_shift_reg_21 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_152, Q => FE_PHN44_spi_com_MISO_shift_21);
  spi_com_MISO_shift_reg_22 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_217, Q => spi_com_MISO_shift(22));
  spi_com_MISO_shift_reg_23 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_219, Q => spi_com_MISO_shift(23));
  spi_com_MISO_shift_reg_24 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_218, Q => FE_PHN23_spi_com_MISO_shift_24);
  spi_com_MISO_shift_reg_25 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_216, Q => spi_com_MISO_shift(25));
  spi_com_MISO_shift_reg_26 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_238, Q => FE_PHN53_spi_com_MISO_shift_26);
  spi_com_MISO_shift_reg_27 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_214, Q => FE_PHN145_spi_com_MISO_shift_27);
  spi_com_MISO_shift_reg_28 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_213, Q => FE_PHN83_spi_com_MISO_shift_28);
  spi_com_MISO_shift_reg_29 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_212, Q => spi_com_MISO_shift(29));
  spi_com_MISO_shift_reg_30 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_210, Q => FE_PHN19_spi_com_MISO_shift_30);
  spi_com_MISO_shift_reg_31 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_209, Q => spi_com_MISO_shift(31));
  spi_com_MISO_shift_reg_32 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_208, Q => spi_com_MISO_shift(32));
  spi_com_MISO_shift_reg_33 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_207, Q => FE_PHN138_spi_com_MISO_shift_33);
  spi_com_MISO_shift_reg_34 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_205, Q => FE_PHN453_spi_com_MISO_shift_34);
  spi_com_MISO_shift_reg_35 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_204, Q => spi_com_MISO_shift(35));
  spi_com_MISO_shift_reg_36 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_202, Q => spi_com_MISO_shift(36));
  spi_com_MISO_shift_reg_37 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_200, Q => FE_PHN11_spi_com_MISO_shift_37);
  spi_com_MISO_shift_reg_38 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_199, Q => FE_PHN25_spi_com_MISO_shift_38);
  spi_com_MISO_shift_reg_39 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_197, Q => FE_PHN152_spi_com_MISO_shift_39);
  spi_com_MISO_shift_reg_40 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_196, Q => spi_com_MISO_shift(40));
  spi_com_MISO_shift_reg_41 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_215, Q => spi_com_MISO_shift(41));
  spi_com_MISO_shift_reg_42 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_236, Q => FE_PHN462_spi_com_MISO_shift_42);
  spi_com_MISO_shift_reg_43 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_194, Q => spi_com_MISO_shift(43));
  spi_com_MISO_shift_reg_44 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_193, Q => FE_PHN155_spi_com_MISO_shift_44);
  spi_com_MISO_shift_reg_45 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_191, Q => spi_com_MISO_shift(45));
  spi_com_MISO_shift_reg_46 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_190, Q => FE_PHN418_spi_com_MISO_shift_46);
  spi_com_MISO_shift_reg_47 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_188, Q => FE_PHN153_spi_com_MISO_shift_47);
  spi_com_MISO_shift_reg_48 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_187, Q => FE_PHN31_spi_com_MISO_shift_48);
  spi_com_MISO_shift_reg_49 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_185, Q => FE_PHN156_spi_com_MISO_shift_49);
  spi_com_MISO_shift_reg_50 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_183, Q => FE_PHN114_spi_com_MISO_shift_50);
  spi_com_MISO_shift_reg_51 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_181, Q => FE_PHN148_spi_com_MISO_shift_51);
  spi_com_MISO_shift_reg_52 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_180, Q => spi_com_MISO_shift(52));
  spi_com_MISO_shift_reg_53 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_179, Q => FE_PHN15_spi_com_MISO_shift_53);
  spi_com_MISO_shift_reg_54 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_177, Q => spi_com_MISO_shift(54));
  spi_com_MISO_shift_reg_55 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_176, Q => FE_PHN87_spi_com_MISO_shift_55);
  spi_com_MISO_shift_reg_56 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_174, Q => spi_com_MISO_shift(56));
  spi_com_MISO_shift_reg_57 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_173, Q => spi_com_MISO_shift(57));
  spi_com_MISO_shift_reg_58 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_195, Q => FE_PHN103_spi_com_MISO_shift_58);
  spi_com_MISO_shift_reg_59 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_169, Q => spi_com_MISO_shift(59));
  spi_com_MISO_shift_reg_60 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_168, Q => FE_PHN42_spi_com_MISO_shift_60);
  spi_com_MISO_shift_reg_61 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_167, Q => FE_PHN115_spi_com_MISO_shift_61);
  spi_com_MISO_shift_reg_62 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_165, Q => spi_com_MISO_shift(62));
  spi_com_MISO_shift_reg_63 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_163, Q => spi_com_MISO_shift(63));
  spi_com_MISO_shift_reg_64 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_162, Q => spi_com_MISO_shift(64));
  spi_com_MISO_shift_reg_65 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_161, Q => FE_PHN102_spi_com_MISO_shift_65);
  spi_com_MISO_shift_reg_66 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_159, Q => FE_PHN16_spi_com_MISO_shift_66);
  spi_com_MISO_shift_reg_67 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_158, Q => spi_com_MISO_shift(67));
  spi_com_MISO_shift_reg_68 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_157, Q => spi_com_MISO_shift(68));
  spi_com_MISO_shift_reg_69 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_155, Q => spi_com_MISO_shift(69));
  spi_com_MISO_shift_reg_70 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_153, Q => FE_PHN21_spi_com_MISO_shift_70);
  spi_com_MISO_shift_reg_71 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_151, Q => spi_com_MISO_shift(71));
  spi_com_MISO_shift_reg_72 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_150, Q => FE_PHN81_spi_com_MISO_shift_72);
  spi_com_MOSI_shift_reg_0 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_186, Q => FE_PHN128_spi_com_MOSI_shift_0);
  spi_com_MOSI_shift_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_234, Q => FE_PHN142_spi_com_MOSI_shift_1);
  spi_com_MOSI_shift_reg_2 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_233, Q => spi_com_MOSI_shift(2));
  spi_com_MOSI_shift_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_232, Q => spi_com_MOSI_shift(3));
  spi_com_MOSI_shift_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_231, Q => spi_com_MOSI_shift(4));
  spi_com_MOSI_shift_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_230, Q => FE_PHN146_spi_com_MOSI_shift_5);
  spi_com_MOSI_shift_reg_6 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_229, Q => spi_com_MOSI_shift(6));
  spi_com_MOSI_shift_reg_7 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_228, Q => FE_PHN131_spi_com_MOSI_shift_7);
  spi_com_MOSI_shift_reg_8 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_242, Q => spi_com_MOSI_shift(8));
  spi_com_MOSI_shift_reg_9 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN302_spi_com_n_226, Q => spi_com_MOSI_shift(9));
  spi_com_MOSI_shift_reg_10 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN294_spi_com_n_247, Q => FE_PHN129_spi_com_MOSI_shift_10);
  spi_com_MOSI_shift_reg_11 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN315_spi_com_n_224, Q => spi_com_MOSI_shift(11));
  spi_com_MOSI_shift_reg_12 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN324_spi_com_n_246, Q => FE_PHN375_spi_com_MOSI_shift_12);
  spi_com_MOSI_shift_reg_13 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_222, Q => spi_com_MOSI_shift(13));
  spi_com_MOSI_shift_reg_14 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_245, Q => FE_PHN379_spi_com_MOSI_shift_14);
  spi_com_SCLK_count_reg_1 : EDFKCND1BWP7T port map(CN => spi_com_n_18, CP => CTS_19, D => FE_PHN371_spi_com_SCLK_count_1, E => FE_PHN229_spi_com_SCLK_count_0, Q => UNCONNECTED0, QN => spi_com_SCLK_count(1));
  spi_com_SCLK_count_reg_2 : DFKCNQD1BWP7T port map(CN => spi_com_n_18, CP => CTS_19, D => FE_PHN292_spi_com_n_43, Q => spi_com_SCLK_count(2));
  spi_com_SCLK_count_reg_3 : DFKCNQD1BWP7T port map(CN => spi_com_n_18, CP => CTS_19, D => FE_PHN303_spi_com_n_55, Q => spi_com_SCLK_count(3));
  spi_com_SCLK_count_reg_4 : DFKCNQD1BWP7T port map(CN => spi_com_n_18, CP => CTS_19, D => FE_PHN288_spi_com_n_129, Q => spi_com_SCLK_count(4));
  spi_com_bit_count_reg_0 : DFXQD1BWP7T port map(CP => CTS_19, DA => spi_com_n_239, DB => spi_com_n_132, Q => spi_com_bit_count(0), SA => FE_PHN419_spi_com_bit_count_0);
  spi_com_bit_count_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN269_spi_com_n_252, Q => spi_com_bit_count(1));
  spi_com_bit_count_reg_3 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN319_spi_com_n_258, Q => spi_com_bit_count(3));
  spi_com_byte_count_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_248, Q => FE_PHN228_spi_com_byte_count_0);
  spi_com_map_data_internal_reg_0 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_116, Q => map_data_volatile(0));
  spi_com_map_data_internal_reg_1 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_115, Q => FE_PHN90_map_data_volatile_1);
  spi_com_map_data_internal_reg_2 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_114, Q => FE_PHN49_map_data_volatile_2);
  spi_com_map_data_internal_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_113, Q => FE_PHN127_map_data_volatile_3);
  spi_com_map_data_internal_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_112, Q => FE_PHN157_map_data_volatile_4);
  spi_com_map_data_internal_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_111, Q => FE_PHN71_map_data_volatile_5);
  spi_com_map_data_internal_reg_6 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_110, Q => map_data_volatile(6));
  spi_com_map_data_internal_reg_7 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_127, Q => map_data_volatile(7));
  spi_com_map_data_internal_reg_8 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_108, Q => FE_PHN124_map_data_volatile_8);
  spi_com_map_data_internal_reg_9 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_107, Q => FE_PHN116_map_data_volatile_9);
  spi_com_map_data_internal_reg_10 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_106, Q => FE_PHN364_map_data_volatile_10);
  spi_com_map_data_internal_reg_11 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_105, Q => FE_PHN125_map_data_volatile_11);
  spi_com_map_data_internal_reg_12 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_104, Q => FE_PHN98_map_data_volatile_12);
  spi_com_map_data_internal_reg_13 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_103, Q => FE_PHN36_map_data_volatile_13);
  spi_com_map_data_internal_reg_14 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_102, Q => FE_PHN55_map_data_volatile_14);
  spi_com_map_data_internal_reg_15 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_100, Q => FE_PHN86_map_data_volatile_15);
  spi_com_map_data_internal_reg_16 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_99, Q => FE_PHN137_map_data_volatile_16);
  spi_com_map_data_internal_reg_17 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_98, Q => map_data_volatile(17));
  spi_com_map_data_internal_reg_18 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_97, Q => FE_PHN77_map_data_volatile_18);
  spi_com_map_data_internal_reg_19 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_96, Q => map_data_volatile(19));
  spi_com_map_data_internal_reg_20 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_95, Q => FE_PHN134_map_data_volatile_20);
  spi_com_map_data_internal_reg_21 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_126, Q => FE_PHN111_map_data_volatile_21);
  spi_com_map_data_internal_reg_22 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_93, Q => FE_PHN110_map_data_volatile_22);
  spi_com_map_data_internal_reg_23 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_92, Q => FE_PHN150_map_data_volatile_23);
  spi_com_map_data_internal_reg_24 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_73, Q => map_data_volatile(24));
  spi_com_map_data_internal_reg_25 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_90, Q => FE_PHN133_map_data_volatile_25);
  spi_com_map_data_internal_reg_26 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_89, Q => map_data_volatile(26));
  spi_com_map_data_internal_reg_27 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_88, Q => map_data_volatile(27));
  spi_com_map_data_internal_reg_28 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_87, Q => map_data_volatile(28));
  spi_com_map_data_internal_reg_29 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_86, Q => FE_PHN59_map_data_volatile_29);
  spi_com_map_data_internal_reg_30 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_85, Q => FE_PHN82_map_data_volatile_30);
  spi_com_map_data_internal_reg_31 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_81, Q => FE_PHN78_map_data_volatile_31);
  spi_com_map_data_internal_reg_32 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_84, Q => FE_PHN106_map_data_volatile_32);
  spi_com_map_data_internal_reg_33 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN405_spi_com_n_83, Q => FE_PHN183_map_data_volatile_33);
  spi_com_map_data_internal_reg_34 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_82, Q => FE_PHN56_map_data_volatile_34);
  spi_com_map_data_internal_reg_35 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_80, Q => FE_PHN147_map_data_volatile_35);
  spi_com_map_data_internal_reg_36 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_79, Q => FE_PHN178_map_data_volatile_36);
  spi_com_map_data_internal_reg_37 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_78, Q => map_data_volatile(37));
  spi_com_map_data_internal_reg_38 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_120, Q => FE_PHN130_map_data_volatile_38);
  spi_com_map_data_internal_reg_39 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_77, Q => FE_PHN119_map_data_volatile_39);
  spi_com_map_data_internal_reg_40 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_76, Q => FE_PHN109_map_data_volatile_40);
  spi_com_map_data_internal_reg_41 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_123, Q => map_data_volatile(41));
  spi_com_map_data_internal_reg_42 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_75, Q => FE_PHN89_map_data_volatile_42);
  spi_com_map_data_internal_reg_43 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_125, Q => FE_PHN108_map_data_volatile_43);
  spi_com_map_data_internal_reg_44 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN494_spi_com_n_74, Q => map_data_volatile(44));
  spi_com_map_data_internal_reg_45 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_91, Q => FE_PHN118_map_data_volatile_45);
  spi_com_map_data_internal_reg_46 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_109, Q => map_data_volatile(46));
  spi_com_map_data_internal_reg_47 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_71, Q => FE_PHN73_map_data_volatile_47);
  spi_com_map_data_internal_reg_48 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_70, Q => FE_PHN50_map_data_volatile_48);
  spi_com_map_data_internal_reg_49 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_69, Q => FE_PHN76_map_data_volatile_49);
  spi_com_map_data_internal_reg_50 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_118, Q => FE_PHN65_map_data_volatile_50);
  spi_com_map_data_internal_reg_51 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN290_spi_com_n_101, Q => map_data_volatile(51));
  spi_com_map_data_internal_reg_52 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_68, Q => FE_PHN154_map_data_volatile_52);
  spi_com_map_data_internal_reg_53 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_67, Q => FE_PHN139_map_data_volatile_53);
  spi_com_map_data_internal_reg_54 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_66, Q => map_data_volatile(54));
  spi_com_map_data_internal_reg_55 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_65, Q => FE_PHN99_map_data_volatile_55);
  spi_com_map_data_internal_reg_56 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_58, Q => map_data_volatile(56));
  spi_com_map_data_internal_reg_57 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_64, Q => FE_PHN132_map_data_volatile_57);
  spi_com_map_data_internal_reg_58 : DFQD1BWP7T port map(CP => CTS_21, D => spi_com_n_72, Q => FE_PHN158_map_data_volatile_58);
  spi_com_map_data_internal_reg_59 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_63, Q => map_data_volatile(59));
  spi_com_map_data_internal_reg_60 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_62, Q => FE_PHN38_map_data_volatile_60);
  spi_com_map_data_internal_reg_61 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_94, Q => FE_PHN104_map_data_volatile_61);
  spi_com_map_data_internal_reg_62 : DFQD1BWP7T port map(CP => CTS_22, D => spi_com_n_61, Q => FE_PHN113_map_data_volatile_62);
  spi_com_map_data_internal_reg_63 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_60, Q => FE_PHN85_map_data_volatile_63);
  spi_com_map_data_internal_reg_64 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_59, Q => map_data_volatile(64));
  spi_com_map_data_internal_reg_65 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_117, Q => map_data_volatile(65));
  spi_com_map_data_internal_reg_66 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_119, Q => map_data_volatile(66));
  spi_com_map_data_internal_reg_67 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_121, Q => map_data_volatile(67));
  spi_com_map_data_internal_reg_68 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_57, Q => FE_PHN48_map_data_volatile_68);
  spi_com_map_data_internal_reg_69 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_56, Q => FE_PHN88_map_data_volatile_69);
  spi_com_map_data_internal_reg_70 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_122, Q => FE_PHN58_map_data_volatile_70);
  spi_com_map_data_internal_reg_71 : DFQD1BWP7T port map(CP => CTS_20, D => spi_com_n_124, Q => FE_PHN177_map_data_volatile_71);
  spi_com_pause_count_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => spi_com_n_244, Q => FE_PHN218_spi_com_pause_count_0);
  spi_com_pause_count_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN260_spi_com_n_255, Q => spi_com_pause_count(1));
  spi_com_state_reg_2 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN334_spi_com_n_45, Q => spi_com_state(2));
  spi_com_g10849 : AO211D0BWP7T port map(A1 => spi_com_n_54, A2 => spi_com_n_141, B => spi_com_n_253, C => spi_com_n_131, Z => spi_com_n_263);
  spi_com_g10850 : IOA21D1BWP7T port map(A1 => spi_com_n_250, A2 => MISO, B => spi_com_n_259, ZN => spi_com_n_262);
  spi_com_g10857 : OAI32D1BWP7T port map(A1 => spi_com_byte_count(2), A2 => spi_com_n_12, A3 => spi_com_n_148, B1 => spi_com_n_2, B2 => spi_com_n_251, ZN => spi_com_n_261);
  spi_com_g10858 : AO21D0BWP7T port map(A1 => spi_com_n_249, A2 => spi_com_bit_count(2), B => spi_com_n_0, Z => spi_com_n_260);
  spi_com_g10859 : IND3D1BWP7T port map(A1 => spi_com_n_250, B1 => spi_com_MISO_shift(0), B2 => spi_com_n_18, ZN => spi_com_n_259);
  spi_com_g10860 : AO22D0BWP7T port map(A1 => spi_com_n_249, A2 => spi_com_bit_count(3), B1 => spi_com_n_46, B2 => spi_com_n_132, Z => spi_com_n_258);
  spi_com_g10861 : OAI22D0BWP7T port map(A1 => spi_com_n_251, A2 => spi_com_n_4, B1 => spi_com_n_148, B2 => spi_com_n_30, ZN => spi_com_n_257);
  spi_com_g10868 : MOAI22D0BWP7T port map(A1 => spi_com_n_133, A2 => spi_com_n_36, B1 => spi_com_n_241, B2 => spi_com_pause_count(2), ZN => spi_com_n_256);
  spi_com_g10869 : IOA21D1BWP7T port map(A1 => spi_com_n_241, A2 => spi_com_pause_count(1), B => spi_com_n_145, ZN => spi_com_n_255);
  spi_com_g10870 : ND3D0BWP7T port map(A1 => spi_com_n_144, A2 => spi_com_n_237, A3 => spi_com_n_135, ZN => spi_com_n_254);
  spi_com_g10871 : NR3D0BWP7T port map(A1 => spi_com_n_240, A2 => spi_com_n_47, A3 => spi_com_n_42, ZN => spi_com_n_253);
  spi_com_g10872 : AO22D0BWP7T port map(A1 => spi_com_n_239, A2 => spi_com_bit_count(1), B1 => spi_com_n_22, B2 => spi_com_n_132, Z => spi_com_n_252);
  spi_com_g10921 : MOAI22D0BWP7T port map(A1 => spi_com_n_148, A2 => spi_com_byte_count(0), B1 => spi_com_n_149, B2 => spi_com_byte_count(0), ZN => spi_com_n_248);
  spi_com_g10922 : ND2D1BWP7T port map(A1 => spi_com_n_225, A2 => spi_com_n_24, ZN => spi_com_n_247);
  spi_com_g10923 : ND2D1BWP7T port map(A1 => spi_com_n_223, A2 => spi_com_n_24, ZN => spi_com_n_246);
  spi_com_g10924 : ND2D1BWP7T port map(A1 => spi_com_n_221, A2 => spi_com_n_24, ZN => spi_com_n_245);
  spi_com_g10925 : IOA21D1BWP7T port map(A1 => spi_com_n_146, A2 => spi_com_pause_count(0), B => spi_com_n_143, ZN => spi_com_n_244);
  spi_com_g10926 : MOAI22D0BWP7T port map(A1 => spi_com_n_148, A2 => spi_com_n_38, B1 => spi_com_n_149, B2 => spi_com_byte_count(1), ZN => FE_PHN306_spi_com_n_243);
  spi_com_g10927 : ND2D1BWP7T port map(A1 => spi_com_n_227, A2 => spi_com_n_24, ZN => FE_PHN301_spi_com_n_242);
  spi_com_g10928 : AOI21D0BWP7T port map(A1 => spi_com_n_147, A2 => spi_com_n_12, B => spi_com_n_149, ZN => spi_com_n_251);
  spi_com_g10929 : AO21D0BWP7T port map(A1 => spi_com_n_54, A2 => spi_com_n_140, B => spi_com_n_240, Z => spi_com_n_250);
  spi_com_g10931 : AO21D0BWP7T port map(A1 => spi_com_n_132, A2 => spi_com_n_19, B => spi_com_n_239, Z => spi_com_n_249);
  spi_com_g10968 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(26), B1 => FE_PHN69_spi_com_MISO_shift_25, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_238);
  spi_com_g10969 : OAI211D1BWP7T port map(A1 => spi_com_n_40, A2 => spi_com_n_136, B => spi_com_n_48, C => spi_com_n_28, ZN => spi_com_n_237);
  spi_com_g10970 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN455_spi_com_MISO_shift_42, B1 => FE_PHN51_spi_com_MISO_shift_41, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_236);
  spi_com_g10971 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(6), B1 => FE_PHN8_spi_com_MISO_shift_5, B2 => spi_com_n_131, Z => spi_com_n_235);
  spi_com_g10972 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(1), B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(0), C1 => spi_com_n_23, C2 => xplayer(1), Z => spi_com_n_234);
  spi_com_g10973 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN75_spi_com_MOSI_shift_2, B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(1), C1 => spi_com_n_23, C2 => xplayer(2), Z => spi_com_n_233);
  spi_com_g10974 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN92_spi_com_MOSI_shift_3, B1 => spi_com_n_131, B2 => FE_PHN75_spi_com_MOSI_shift_2, C1 => spi_com_n_23, C2 => xplayer(3), Z => spi_com_n_232);
  spi_com_g10975 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN96_spi_com_MOSI_shift_4, B1 => spi_com_n_131, B2 => FE_PHN92_spi_com_MOSI_shift_3, C1 => spi_com_n_23, C2 => yplayer(0), Z => spi_com_n_231);
  spi_com_g10976 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(5), B1 => spi_com_n_131, B2 => FE_PHN96_spi_com_MOSI_shift_4, C1 => spi_com_n_23, C2 => yplayer(1), Z => spi_com_n_230);
  spi_com_g10977 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN112_spi_com_MOSI_shift_6, B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(5), C1 => spi_com_n_23, C2 => yplayer(2), Z => FE_PHN295_spi_com_n_229);
  spi_com_g10978 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(7), B1 => spi_com_n_131, B2 => FE_PHN112_spi_com_MOSI_shift_6, C1 => spi_com_n_23, C2 => yplayer(3), Z => spi_com_n_228);
  spi_com_g10979 : AOI222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(8), B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(7), C1 => spi_com_n_23, C2 => level_abs(0), ZN => spi_com_n_227);
  spi_com_g10980 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(9), B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(8), C1 => spi_com_n_23, C2 => level_abs(1), Z => spi_com_n_226);
  spi_com_g10981 : AOI222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(10), B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(9), C1 => spi_com_n_23, C2 => level_abs(2), ZN => spi_com_n_225);
  spi_com_g10982 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(11), B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(10), C1 => spi_com_n_23, C2 => level_abs(3), Z => spi_com_n_224);
  spi_com_g10983 : AOI222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(12), B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(11), C1 => spi_com_n_23, C2 => level_abs(4), ZN => spi_com_n_223);
  spi_com_g10984 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN141_spi_com_MOSI_shift_13, B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(12), C1 => MOSI_data(13), C2 => spi_com_n_23, Z => spi_com_n_222);
  spi_com_g10985 : AOI222D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(14), B1 => spi_com_n_131, B2 => FE_PHN141_spi_com_MOSI_shift_13, C1 => dir_mined(0), C2 => spi_com_n_23, ZN => spi_com_n_221);
  spi_com_g10986 : AO222D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN175_spi_com_n_9, B1 => spi_com_n_131, B2 => spi_com_MOSI_shift(14), C1 => dir_mined(1), C2 => spi_com_n_23, Z => spi_com_n_220);
  spi_com_g10987 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN27_spi_com_MISO_shift_23, B1 => FE_PHN35_spi_com_MISO_shift_22, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_219);
  spi_com_g10988 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(24), B1 => FE_PHN27_spi_com_MISO_shift_23, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_218);
  spi_com_g10989 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN35_spi_com_MISO_shift_22, B1 => spi_com_MISO_shift(21), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_217);
  spi_com_g10990 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN69_spi_com_MISO_shift_25, B1 => spi_com_MISO_shift(24), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_216);
  spi_com_g10991 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN51_spi_com_MISO_shift_41, B1 => FE_PHN170_spi_com_MISO_shift_40, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_215);
  spi_com_g10992 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(27), B1 => spi_com_MISO_shift(26), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_214);
  spi_com_g10993 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(28), B1 => spi_com_MISO_shift(27), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_213);
  spi_com_g10994 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN40_spi_com_MISO_shift_29, B1 => spi_com_MISO_shift(28), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_212);
  spi_com_g10995 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(1), B1 => spi_com_MISO_shift(0), B2 => spi_com_n_131, Z => spi_com_n_211);
  spi_com_g10996 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(30), B1 => FE_PHN40_spi_com_MISO_shift_29, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_210);
  spi_com_g10997 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN29_spi_com_MISO_shift_31, B1 => spi_com_MISO_shift(30), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_209);
  spi_com_g10998 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN62_spi_com_MISO_shift_32, B1 => FE_PHN29_spi_com_MISO_shift_31, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_208);
  spi_com_g10999 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(33), B1 => FE_PHN62_spi_com_MISO_shift_32, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_207);
  spi_com_g11000 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(2), B1 => spi_com_MISO_shift(1), B2 => spi_com_n_131, Z => spi_com_n_206);
  spi_com_g11001 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(34), B1 => spi_com_MISO_shift(33), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_205);
  spi_com_g11002 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN57_spi_com_MISO_shift_35, B1 => spi_com_MISO_shift(34), B2 => spi_com_n_131, Z => spi_com_n_204);
  spi_com_g11003 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(3), B1 => spi_com_MISO_shift(2), B2 => spi_com_n_131, Z => spi_com_n_203);
  spi_com_g11004 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN20_spi_com_MISO_shift_36, B1 => FE_PHN57_spi_com_MISO_shift_35, B2 => spi_com_n_131, Z => spi_com_n_202);
  spi_com_g11005 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(4), B1 => spi_com_MISO_shift(3), B2 => spi_com_n_131, Z => spi_com_n_201);
  spi_com_g11006 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(37), B1 => FE_PHN20_spi_com_MISO_shift_36, B2 => spi_com_n_131, Z => spi_com_n_200);
  spi_com_g11007 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(38), B1 => spi_com_MISO_shift(37), B2 => spi_com_n_131, Z => spi_com_n_199);
  spi_com_g11008 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN8_spi_com_MISO_shift_5, B1 => spi_com_MISO_shift(4), B2 => spi_com_n_131, Z => spi_com_n_198);
  spi_com_g11009 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(39), B1 => spi_com_MISO_shift(38), B2 => spi_com_n_131, Z => spi_com_n_197);
  spi_com_g11010 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN170_spi_com_MISO_shift_40, B1 => spi_com_MISO_shift(39), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_196);
  spi_com_g11011 : IND2D1BWP7T port map(A1 => spi_com_n_146, B1 => spi_com_n_143, ZN => spi_com_n_241);
  spi_com_g11012 : NR3D0BWP7T port map(A1 => spi_com_n_141, A2 => spi_com_n_40, A3 => spi_com_n_34, ZN => spi_com_n_240);
  spi_com_g11013 : AOI211XD0BWP7T port map(A1 => spi_com_n_138, A2 => spi_com_n_26, B => spi_com_n_132, C => spi_com_n_17, ZN => spi_com_n_239);
  spi_com_g11014 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(58), B1 => FE_PHN107_spi_com_MISO_shift_57, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_195);
  spi_com_g11015 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN54_spi_com_MISO_shift_43, B1 => spi_com_MISO_shift(42), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_194);
  spi_com_g11016 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(44), B1 => FE_PHN54_spi_com_MISO_shift_43, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_193);
  spi_com_g11017 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN12_spi_com_MISO_shift_8, B1 => spi_com_MISO_shift(7), B2 => spi_com_n_131, Z => spi_com_n_192);
  spi_com_g11018 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN67_spi_com_MISO_shift_45, B1 => spi_com_MISO_shift(44), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_191);
  spi_com_g11019 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(46), B1 => FE_PHN67_spi_com_MISO_shift_45, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_190);
  spi_com_g11020 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(9), B1 => FE_PHN12_spi_com_MISO_shift_8, B2 => spi_com_n_131, Z => spi_com_n_189);
  spi_com_g11021 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(47), B1 => spi_com_MISO_shift(46), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_188);
  spi_com_g11022 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(48), B1 => spi_com_MISO_shift(47), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_187);
  spi_com_g11023 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MOSI_shift(0), B1 => xplayer(0), B2 => spi_com_n_23, Z => spi_com_n_186);
  spi_com_g11024 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(49), B1 => spi_com_MISO_shift(48), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_185);
  spi_com_g11025 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(10), B1 => spi_com_MISO_shift(9), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_184);
  spi_com_g11026 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(50), B1 => spi_com_MISO_shift(49), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_183);
  spi_com_g11027 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(11), B1 => spi_com_MISO_shift(10), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_182);
  spi_com_g11028 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(51), B1 => spi_com_MISO_shift(50), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_181);
  spi_com_g11029 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN117_spi_com_MISO_shift_52, B1 => spi_com_MISO_shift(51), B2 => spi_com_n_131, Z => spi_com_n_180);
  spi_com_g11030 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(53), B1 => FE_PHN117_spi_com_MISO_shift_52, B2 => spi_com_n_131, Z => spi_com_n_179);
  spi_com_g11031 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN187_spi_com_MISO_shift_12, B1 => spi_com_MISO_shift(11), B2 => FE_OFN6_spi_com_n_131, Z => FE_PHN406_spi_com_n_178);
  spi_com_g11032 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN37_spi_com_MISO_shift_54, B1 => spi_com_MISO_shift(53), B2 => spi_com_n_131, Z => spi_com_n_177);
  spi_com_g11033 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(55), B1 => FE_PHN37_spi_com_MISO_shift_54, B2 => spi_com_n_131, Z => spi_com_n_176);
  spi_com_g11034 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(13), B1 => FE_PHN187_spi_com_MISO_shift_12, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_175);
  spi_com_g11035 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN14_spi_com_MISO_shift_56, B1 => spi_com_MISO_shift(55), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_174);
  spi_com_g11036 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN107_spi_com_MISO_shift_57, B1 => FE_PHN14_spi_com_MISO_shift_56, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_173);
  spi_com_g11037 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(7), B1 => spi_com_MISO_shift(6), B2 => spi_com_n_131, Z => spi_com_n_172);
  spi_com_g11038 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN441_spi_com_MISO_shift_14, B1 => spi_com_MISO_shift(13), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_171);
  spi_com_g11039 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN30_spi_com_MISO_shift_15, B1 => FE_PHN190_spi_com_MISO_shift_14, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_170);
  spi_com_g11040 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN26_spi_com_MISO_shift_59, B1 => spi_com_MISO_shift(58), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_169);
  spi_com_g11041 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(60), B1 => FE_PHN26_spi_com_MISO_shift_59, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_168);
  spi_com_g11042 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(61), B1 => spi_com_MISO_shift(60), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_167);
  spi_com_g11043 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN10_spi_com_MISO_shift_16, B1 => FE_PHN30_spi_com_MISO_shift_15, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_166);
  spi_com_g11044 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN149_spi_com_MISO_shift_62, B1 => spi_com_MISO_shift(61), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_165);
  spi_com_g11045 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(17), B1 => FE_PHN10_spi_com_MISO_shift_16, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_164);
  spi_com_g11046 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN9_spi_com_MISO_shift_63, B1 => FE_PHN149_spi_com_MISO_shift_62, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_163);
  spi_com_g11047 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN151_spi_com_MISO_shift_64, B1 => FE_PHN9_spi_com_MISO_shift_63, B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_162);
  spi_com_g11048 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(65), B1 => FE_PHN151_spi_com_MISO_shift_64, B2 => spi_com_n_131, Z => spi_com_n_161);
  spi_com_g11049 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => FE_PHN398_spi_com_MISO_shift_18, B1 => spi_com_MISO_shift(17), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_160);
  spi_com_g11050 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(66), B1 => spi_com_MISO_shift(65), B2 => spi_com_n_131, Z => spi_com_n_159);
  spi_com_g11051 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN32_spi_com_MISO_shift_67, B1 => spi_com_MISO_shift(66), B2 => spi_com_n_131, Z => spi_com_n_158);
  spi_com_g11052 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN28_spi_com_MISO_shift_68, B1 => FE_PHN32_spi_com_MISO_shift_67, B2 => spi_com_n_131, Z => spi_com_n_157);
  spi_com_g11053 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(19), B1 => spi_com_MISO_shift(18), B2 => spi_com_n_131, Z => spi_com_n_156);
  spi_com_g11054 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN13_spi_com_MISO_shift_69, B1 => FE_PHN28_spi_com_MISO_shift_68, B2 => spi_com_n_131, Z => spi_com_n_155);
  spi_com_g11055 : AO22D0BWP7T port map(A1 => FE_OFN5_spi_com_n_139, A2 => spi_com_MISO_shift(20), B1 => spi_com_MISO_shift(19), B2 => FE_OFN6_spi_com_n_131, Z => spi_com_n_154);
  spi_com_g11056 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(70), B1 => FE_PHN13_spi_com_MISO_shift_69, B2 => spi_com_n_131, Z => spi_com_n_153);
  spi_com_g11057 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(21), B1 => spi_com_MISO_shift(20), B2 => spi_com_n_131, Z => spi_com_n_152);
  spi_com_g11058 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => FE_PHN24_spi_com_MISO_shift_71, B1 => spi_com_MISO_shift(70), B2 => spi_com_n_131, Z => spi_com_n_151);
  spi_com_g11059 : AO22D0BWP7T port map(A1 => spi_com_n_139, A2 => spi_com_MISO_shift(72), B1 => FE_PHN24_spi_com_MISO_shift_71, B2 => spi_com_n_131, Z => spi_com_n_150);
  spi_com_g11060 : INVD1BWP7T port map(I => spi_com_n_147, ZN => spi_com_n_148);
  spi_com_g11061 : NR2D1BWP7T port map(A1 => spi_com_n_142, A2 => spi_com_n_17, ZN => spi_com_n_149);
  spi_com_g11062 : INR2XD0BWP7T port map(A1 => spi_com_n_142, B1 => spi_com_n_49, ZN => spi_com_n_147);
  spi_com_g11063 : IND3D1BWP7T port map(A1 => spi_com_pause_count(1), B1 => spi_com_pause_count(0), B2 => spi_com_n_134, ZN => spi_com_n_145);
  spi_com_g11064 : AOI22D0BWP7T port map(A1 => spi_com_n_54, A2 => spi_com_n_130, B1 => spi_com_n_137, B2 => spi_com_n_27, ZN => spi_com_n_144);
  spi_com_g11065 : OAI211D1BWP7T port map(A1 => spi_com_n_28, A2 => spi_com_n_130, B => spi_com_n_13, C => spi_com_n_25, ZN => spi_com_n_146);
  spi_com_g11066 : IND2D1BWP7T port map(A1 => spi_com_pause_count(0), B1 => spi_com_n_134, ZN => spi_com_n_143);
  spi_com_g11067 : NR2XD0BWP7T port map(A1 => spi_com_n_137, A2 => spi_com_n_28, ZN => spi_com_n_142);
  spi_com_g11069 : INVD1BWP7T port map(I => spi_com_n_140, ZN => spi_com_n_141);
  spi_com_g11071 : NR2XD0BWP7T port map(A1 => spi_com_n_138, A2 => spi_com_n_128, ZN => spi_com_n_140);
  spi_com_g11072 : ND2D1P5BWP7T port map(A1 => spi_com_n_135, A2 => spi_com_n_14, ZN => spi_com_n_139);
  spi_com_g11073 : NR2XD0BWP7T port map(A1 => spi_com_n_128, A2 => spi_com_n_34, ZN => spi_com_n_136);
  spi_com_g11074 : INR2XD0BWP7T port map(A1 => spi_com_n_35, B1 => spi_com_n_128, ZN => spi_com_n_138);
  spi_com_g11075 : ND2D1BWP7T port map(A1 => spi_com_n_130, A2 => spi_com_n_29, ZN => spi_com_n_137);
  spi_com_g11076 : INVD0BWP7T port map(I => spi_com_n_134, ZN => spi_com_n_133);
  spi_com_g11078 : IND2D1BWP7T port map(A1 => spi_com_n_13, B1 => spi_com_n_128, ZN => spi_com_n_135);
  spi_com_g11079 : NR3D0BWP7T port map(A1 => spi_com_n_128, A2 => spi_com_n_29, A3 => spi_com_n_28, ZN => spi_com_n_134);
  spi_com_g11080 : NR3D0BWP7T port map(A1 => spi_com_n_128, A2 => spi_com_n_35, A3 => spi_com_n_25, ZN => spi_com_n_132);
  spi_com_g11081 : NR2XD1BWP7T port map(A1 => spi_com_n_128, A2 => spi_com_n_13, ZN => spi_com_n_131);
  spi_com_g11082 : INVD1BWP7T port map(I => spi_com_n_128, ZN => spi_com_n_130);
  spi_com_g11084 : MOAI22D0BWP7T port map(A1 => spi_com_n_53, A2 => spi_com_SCLK_count(4), B1 => spi_com_n_53, B2 => spi_com_SCLK_count(4), ZN => spi_com_n_129);
  spi_com_g11157 : IND2D1BWP7T port map(A1 => spi_com_n_53, B1 => spi_com_SCLK_count(4), ZN => spi_com_n_128);
  spi_com_g11158 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN52_map_data_volatile_7, B1 => FE_PHN12_spi_com_MISO_shift_8, B2 => spi_com_n_51, Z => spi_com_n_127);
  spi_com_g11159 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(21), B1 => FE_PHN35_spi_com_MISO_shift_22, B2 => spi_com_n_51, Z => spi_com_n_126);
  spi_com_g11160 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(43), B1 => spi_com_MISO_shift(44), B2 => spi_com_n_51, Z => spi_com_n_125);
  spi_com_g11161 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN385_map_data_volatile_71, B1 => spi_com_MISO_shift(72), B2 => spi_com_n_51, Z => spi_com_n_124);
  spi_com_g11162 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN122_map_data_volatile_41, B1 => FE_PHN455_spi_com_MISO_shift_42, B2 => spi_com_n_51, Z => spi_com_n_123);
  spi_com_g11163 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(70), B1 => FE_PHN24_spi_com_MISO_shift_71, B2 => spi_com_n_51, Z => spi_com_n_122);
  spi_com_g11164 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN60_map_data_volatile_67, B1 => FE_PHN28_spi_com_MISO_shift_68, B2 => spi_com_n_51, Z => spi_com_n_121);
  spi_com_g11165 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(38), B1 => spi_com_MISO_shift(39), B2 => spi_com_n_51, Z => spi_com_n_120);
  spi_com_g11166 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN70_map_data_volatile_66, B1 => FE_PHN32_spi_com_MISO_shift_67, B2 => spi_com_n_51, Z => spi_com_n_119);
  spi_com_g11167 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(50), B1 => spi_com_MISO_shift(51), B2 => spi_com_n_51, Z => spi_com_n_118);
  spi_com_g11168 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN33_map_data_volatile_65, B1 => spi_com_MISO_shift(66), B2 => spi_com_n_51, Z => spi_com_n_117);
  spi_com_g11169 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN95_map_data_volatile_0, B1 => spi_com_MISO_shift(1), B2 => spi_com_n_51, Z => spi_com_n_116);
  spi_com_g11170 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(1), B1 => spi_com_MISO_shift(2), B2 => spi_com_n_51, Z => spi_com_n_115);
  spi_com_g11171 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(2), B1 => spi_com_MISO_shift(3), B2 => spi_com_n_51, Z => spi_com_n_114);
  spi_com_g11172 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(3), B1 => spi_com_MISO_shift(4), B2 => spi_com_n_51, Z => spi_com_n_113);
  spi_com_g11173 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(4), B1 => FE_PHN8_spi_com_MISO_shift_5, B2 => spi_com_n_51, Z => spi_com_n_112);
  spi_com_g11174 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(5), B1 => spi_com_MISO_shift(6), B2 => spi_com_n_51, Z => spi_com_n_111);
  spi_com_g11175 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN94_map_data_volatile_6, B1 => spi_com_MISO_shift(7), B2 => spi_com_n_51, Z => spi_com_n_110);
  spi_com_g11176 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN381_map_data_volatile_46, B1 => spi_com_MISO_shift(47), B2 => spi_com_n_51, Z => spi_com_n_109);
  spi_com_g11177 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(8), B1 => spi_com_MISO_shift(9), B2 => spi_com_n_51, Z => spi_com_n_108);
  spi_com_g11178 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(9), B1 => spi_com_MISO_shift(10), B2 => spi_com_n_51, Z => spi_com_n_107);
  spi_com_g11179 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(10), B1 => FE_PHN409_spi_com_MISO_shift_11, B2 => spi_com_n_51, Z => spi_com_n_106);
  spi_com_g11180 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(11), B1 => FE_PHN187_spi_com_MISO_shift_12, B2 => spi_com_n_51, Z => spi_com_n_105);
  spi_com_g11181 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(12), B1 => spi_com_MISO_shift(13), B2 => spi_com_n_51, Z => spi_com_n_104);
  spi_com_g11182 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(13), B1 => FE_PHN190_spi_com_MISO_shift_14, B2 => spi_com_n_51, Z => spi_com_n_103);
  spi_com_g11183 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(14), B1 => FE_PHN30_spi_com_MISO_shift_15, B2 => spi_com_n_51, Z => spi_com_n_102);
  spi_com_g11184 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(51), B1 => FE_PHN117_spi_com_MISO_shift_52, B2 => spi_com_n_51, Z => spi_com_n_101);
  spi_com_g11185 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(15), B1 => FE_PHN10_spi_com_MISO_shift_16, B2 => spi_com_n_51, Z => spi_com_n_100);
  spi_com_g11186 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(16), B1 => spi_com_MISO_shift(17), B2 => spi_com_n_51, Z => spi_com_n_99);
  spi_com_g11187 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN61_map_data_volatile_17, B1 => FE_PHN398_spi_com_MISO_shift_18, B2 => spi_com_n_51, Z => spi_com_n_98);
  spi_com_g11188 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(18), B1 => spi_com_MISO_shift(19), B2 => spi_com_n_51, Z => spi_com_n_97);
  spi_com_g11189 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN43_map_data_volatile_19, B1 => spi_com_MISO_shift(20), B2 => spi_com_n_51, Z => spi_com_n_96);
  spi_com_g11190 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(20), B1 => spi_com_MISO_shift(21), B2 => spi_com_n_51, Z => spi_com_n_95);
  spi_com_g11191 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(61), B1 => FE_PHN149_spi_com_MISO_shift_62, B2 => spi_com_n_51, Z => spi_com_n_94);
  spi_com_g11192 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(22), B1 => FE_PHN27_spi_com_MISO_shift_23, B2 => spi_com_n_51, Z => spi_com_n_93);
  spi_com_g11193 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(23), B1 => spi_com_MISO_shift(24), B2 => spi_com_n_51, Z => spi_com_n_92);
  spi_com_g11194 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(45), B1 => spi_com_MISO_shift(46), B2 => spi_com_n_51, Z => spi_com_n_91);
  spi_com_g11195 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(25), B1 => spi_com_MISO_shift(26), B2 => spi_com_n_51, Z => spi_com_n_90);
  spi_com_g11196 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN63_map_data_volatile_26, B1 => spi_com_MISO_shift(27), B2 => spi_com_n_51, Z => spi_com_n_89);
  spi_com_g11197 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN41_map_data_volatile_27, B1 => spi_com_MISO_shift(28), B2 => spi_com_n_51, Z => spi_com_n_88);
  spi_com_g11198 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN47_map_data_volatile_28, B1 => FE_PHN40_spi_com_MISO_shift_29, B2 => spi_com_n_51, Z => spi_com_n_87);
  spi_com_g11199 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(29), B1 => spi_com_MISO_shift(30), B2 => spi_com_n_51, Z => spi_com_n_86);
  spi_com_g11200 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(30), B1 => FE_PHN29_spi_com_MISO_shift_31, B2 => spi_com_n_51, Z => spi_com_n_85);
  spi_com_g11201 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(32), B1 => spi_com_MISO_shift(33), B2 => spi_com_n_51, Z => spi_com_n_84);
  spi_com_g11202 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(33), B1 => spi_com_MISO_shift(34), B2 => spi_com_n_51, Z => spi_com_n_83);
  spi_com_g11203 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(34), B1 => FE_PHN57_spi_com_MISO_shift_35, B2 => spi_com_n_51, Z => spi_com_n_82);
  spi_com_g11204 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(31), B1 => FE_PHN62_spi_com_MISO_shift_32, B2 => spi_com_n_51, Z => spi_com_n_81);
  spi_com_g11205 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(35), B1 => FE_PHN20_spi_com_MISO_shift_36, B2 => spi_com_n_51, Z => spi_com_n_80);
  spi_com_g11206 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN377_map_data_volatile_36, B1 => spi_com_MISO_shift(37), B2 => spi_com_n_51, Z => spi_com_n_79);
  spi_com_g11207 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN378_map_data_volatile_37, B1 => spi_com_MISO_shift(38), B2 => spi_com_n_51, Z => spi_com_n_78);
  spi_com_g11208 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(39), B1 => FE_PHN170_spi_com_MISO_shift_40, B2 => spi_com_n_51, Z => spi_com_n_77);
  spi_com_g11209 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(40), B1 => FE_PHN51_spi_com_MISO_shift_41, B2 => spi_com_n_51, Z => spi_com_n_76);
  spi_com_g11210 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(42), B1 => FE_PHN54_spi_com_MISO_shift_43, B2 => spi_com_n_51, Z => spi_com_n_75);
  spi_com_g11211 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(44), B1 => FE_PHN67_spi_com_MISO_shift_45, B2 => spi_com_n_51, Z => spi_com_n_74);
  spi_com_g11212 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN74_map_data_volatile_24, B1 => FE_PHN69_spi_com_MISO_shift_25, B2 => spi_com_n_51, Z => spi_com_n_73);
  spi_com_g11213 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(58), B1 => FE_PHN26_spi_com_MISO_shift_59, B2 => spi_com_n_51, Z => spi_com_n_72);
  spi_com_g11214 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(47), B1 => spi_com_MISO_shift(48), B2 => spi_com_n_51, Z => spi_com_n_71);
  spi_com_g11215 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(48), B1 => spi_com_MISO_shift(49), B2 => spi_com_n_51, Z => spi_com_n_70);
  spi_com_g11216 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(49), B1 => spi_com_MISO_shift(50), B2 => spi_com_n_51, Z => spi_com_n_69);
  spi_com_g11217 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(52), B1 => spi_com_MISO_shift(53), B2 => spi_com_n_51, Z => spi_com_n_68);
  spi_com_g11218 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(53), B1 => FE_PHN37_spi_com_MISO_shift_54, B2 => spi_com_n_51, Z => spi_com_n_67);
  spi_com_g11219 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN84_map_data_volatile_54, B1 => spi_com_MISO_shift(55), B2 => spi_com_n_51, Z => spi_com_n_66);
  spi_com_g11220 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(55), B1 => FE_PHN14_spi_com_MISO_shift_56, B2 => spi_com_n_51, Z => spi_com_n_65);
  spi_com_g11221 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(57), B1 => spi_com_MISO_shift(58), B2 => spi_com_n_51, Z => spi_com_n_64);
  spi_com_g11222 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN45_map_data_volatile_59, B1 => spi_com_MISO_shift(60), B2 => spi_com_n_51, Z => spi_com_n_63);
  spi_com_g11223 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(60), B1 => spi_com_MISO_shift(61), B2 => spi_com_n_51, Z => spi_com_n_62);
  spi_com_g11224 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(62), B1 => FE_PHN9_spi_com_MISO_shift_63, B2 => spi_com_n_51, Z => spi_com_n_61);
  spi_com_g11225 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(63), B1 => FE_PHN151_spi_com_MISO_shift_64, B2 => spi_com_n_51, Z => spi_com_n_60);
  spi_com_g11226 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN39_map_data_volatile_64, B1 => spi_com_MISO_shift(65), B2 => spi_com_n_51, Z => spi_com_n_59);
  spi_com_g11227 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => FE_PHN126_map_data_volatile_56, B1 => FE_PHN107_spi_com_MISO_shift_57, B2 => spi_com_n_51, Z => spi_com_n_58);
  spi_com_g11228 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(68), B1 => FE_PHN13_spi_com_MISO_shift_69, B2 => spi_com_n_51, Z => spi_com_n_57);
  spi_com_g11229 : AO22D0BWP7T port map(A1 => spi_com_n_52, A2 => map_data_volatile(69), B1 => spi_com_MISO_shift(70), B2 => spi_com_n_51, Z => spi_com_n_56);
  spi_com_g11231 : MOAI22D0BWP7T port map(A1 => spi_com_n_41, A2 => spi_com_SCLK_count(3), B1 => spi_com_n_41, B2 => spi_com_SCLK_count(3), ZN => spi_com_n_55);
  spi_com_g11232 : NR2D1BWP7T port map(A1 => spi_com_n_49, A2 => spi_com_n_39, ZN => spi_com_n_54);
  spi_com_g11233 : IND2D1BWP7T port map(A1 => spi_com_n_41, B1 => spi_com_SCLK_count(3), ZN => spi_com_n_53);
  spi_com_g11234 : ND2D2BWP7T port map(A1 => spi_com_n_50, A2 => spi_com_n_32, ZN => spi_com_n_52);
  spi_com_g11235 : IND2D1BWP7T port map(A1 => spi_com_n_39, B1 => spi_com_n_44, ZN => spi_com_n_50);
  spi_com_g11237 : NR2D4BWP7T port map(A1 => spi_com_n_39, A2 => spi_com_n_44, ZN => spi_com_n_51);
  spi_com_g11238 : INVD0BWP7T port map(I => spi_com_n_47, ZN => spi_com_n_48);
  spi_com_g11239 : OAI31D0BWP7T port map(A1 => spi_com_bit_count(3), A2 => spi_com_n_6, A3 => spi_com_n_19, B => spi_com_n_16, ZN => spi_com_n_46);
  spi_com_g11240 : OAI21D0BWP7T port map(A1 => MOSI_data(13), A2 => spi_com_n_33, B => spi_com_n_44, ZN => spi_com_n_49);
  spi_com_g11241 : IND4D0BWP7T port map(A1 => FE_OFN0_reset, B1 => spi_com_n_13, B2 => spi_com_n_39, B3 => spi_com_n_31, ZN => spi_com_n_47);
  spi_com_g11242 : NR2XD0BWP7T port map(A1 => spi_com_n_42, A2 => spi_com_n_20, ZN => spi_com_n_45);
  spi_com_g11244 : MOAI22D0BWP7T port map(A1 => spi_com_n_15, A2 => spi_com_SCLK_count(2), B1 => spi_com_n_15, B2 => spi_com_SCLK_count(2), ZN => spi_com_n_43);
  spi_com_g11245 : ND3D0BWP7T port map(A1 => spi_com_n_37, A2 => spi_com_byte_count(2), A3 => spi_com_byte_count(3), ZN => spi_com_n_44);
  spi_com_g11246 : NR2XD0BWP7T port map(A1 => spi_com_n_40, A2 => spi_com_n_33, ZN => spi_com_n_42);
  spi_com_g11247 : IND2D1BWP7T port map(A1 => spi_com_n_15, B1 => spi_com_SCLK_count(2), ZN => spi_com_n_41);
  spi_com_g11248 : HA1D0BWP7T port map(A => spi_com_byte_count(0), B => spi_com_n_7, CO => spi_com_n_37, S => spi_com_n_38);
  spi_com_g11249 : AOI31D0BWP7T port map(A1 => spi_com_n_8, A2 => spi_com_pause_count(1), A3 => spi_com_pause_count(0), B => spi_com_n_21, ZN => spi_com_n_36);
  spi_com_g11250 : ND2D1BWP7T port map(A1 => spi_com_n_26, A2 => FE_PHN237_spi_com_state_2, ZN => spi_com_n_40);
  spi_com_g11252 : IND2D1BWP7T port map(A1 => FE_PHN237_spi_com_state_2, B1 => spi_com_n_26, ZN => spi_com_n_39);
  spi_com_g11253 : INVD1BWP7T port map(I => spi_com_n_34, ZN => spi_com_n_33);
  spi_com_g11254 : OAI31D0BWP7T port map(A1 => FE_PHN237_spi_com_state_2, A2 => spi_com_state(1), A3 => spi_com_n_3, B => FE_DBTN0_reset, ZN => spi_com_n_32);
  spi_com_g11255 : OAI21D0BWP7T port map(A1 => spi_com_n_10, A2 => spi_com_send_in1, B => spi_com_n_23, ZN => spi_com_n_31);
  spi_com_g11256 : OA32D1BWP7T port map(A1 => spi_com_byte_count(3), A2 => spi_com_n_2, A3 => spi_com_n_12, B1 => spi_com_byte_count(2), B2 => spi_com_n_4, Z => spi_com_n_30);
  spi_com_g11257 : NR3D0BWP7T port map(A1 => spi_com_n_16, A2 => spi_com_bit_count(1), A3 => FE_PHN226_spi_com_bit_count_0, ZN => spi_com_n_35);
  spi_com_g11258 : NR3D0BWP7T port map(A1 => spi_com_n_12, A2 => spi_com_byte_count(2), A3 => spi_com_byte_count(3), ZN => spi_com_n_34);
  spi_com_g11259 : INVD0BWP7T port map(I => spi_com_n_28, ZN => spi_com_n_27);
  spi_com_g11260 : INVD0BWP7T port map(I => spi_com_n_26, ZN => spi_com_n_25);
  spi_com_g11261 : INR2XD0BWP7T port map(A1 => spi_com_n_21, B1 => spi_com_pause_count(0), ZN => spi_com_n_29);
  spi_com_g11262 : IND2D1BWP7T port map(A1 => spi_com_n_14, B1 => spi_com_state(1), ZN => spi_com_n_28);
  spi_com_g11263 : NR2XD0BWP7T port map(A1 => spi_com_n_14, A2 => spi_com_state(1), ZN => spi_com_n_26);
  spi_com_g11264 : CKXOR2D0BWP7T port map(A1 => spi_com_bit_count(1), A2 => FE_PHN226_spi_com_bit_count_0, Z => spi_com_n_22);
  spi_com_g11265 : ND3D0BWP7T port map(A1 => SS, A2 => FE_PHN237_spi_com_state_2, A3 => FE_DBTN0_reset, ZN => spi_com_n_24);
  spi_com_g11266 : CKAN2D1BWP7T port map(A1 => SS, A2 => spi_com_n_20, Z => spi_com_n_23);
  spi_com_g11267 : INVD0BWP7T port map(I => spi_com_n_18, ZN => spi_com_n_17);
  spi_com_g11268 : NR2XD0BWP7T port map(A1 => spi_com_n_8, A2 => spi_com_pause_count(1), ZN => spi_com_n_21);
  spi_com_g11269 : NR2XD0BWP7T port map(A1 => FE_PHN237_spi_com_state_2, A2 => FE_OFN0_reset, ZN => spi_com_n_20);
  spi_com_g11270 : ND2D1BWP7T port map(A1 => spi_com_bit_count(1), A2 => FE_PHN226_spi_com_bit_count_0, ZN => spi_com_n_19);
  spi_com_g11271 : NR2XD0BWP7T port map(A1 => SS, A2 => FE_OFN0_reset, ZN => spi_com_n_18);
  spi_com_g11272 : CKND2D1BWP7T port map(A1 => spi_com_n_6, A2 => spi_com_bit_count(3), ZN => spi_com_n_16);
  spi_com_g11273 : IND2D1BWP7T port map(A1 => FE_PHN240_spi_com_SCLK_count_1, B1 => FE_PHN229_spi_com_SCLK_count_0, ZN => spi_com_n_15);
  spi_com_g11274 : ND2D1BWP7T port map(A1 => spi_com_state(0), A2 => FE_DBTN0_reset, ZN => spi_com_n_14);
  spi_com_g11275 : ND2D1BWP7T port map(A1 => SCLK, A2 => FE_DBTN0_reset, ZN => spi_com_n_13);
  spi_com_g11276 : ND2D1BWP7T port map(A1 => spi_com_byte_count(1), A2 => spi_com_byte_count(0), ZN => spi_com_n_12);
  spi_com_MOSI_shift_reg_15 : DFD0BWP7T port map(CP => CTS_19, D => spi_com_n_220, Q => spi_com_n_9, QN => spi_com_n_1);
  spi_com_SCLK_count_reg_0 : DFKCND1BWP7T port map(CN => spi_com_n_5, CP => CTS_19, D => spi_com_n_18, Q => spi_com_SCLK_count(0), QN => FE_PHN180_spi_com_n_5);
  spi_com_bit_count_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN275_spi_com_n_260, Q => spi_com_bit_count(2), QN => spi_com_n_6);
  spi_com_byte_count_reg_1 : DFD1BWP7T port map(CP => CTS_19, D => spi_com_n_243, Q => spi_com_byte_count(1), QN => spi_com_n_7);
  spi_com_byte_count_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN256_spi_com_n_261, Q => spi_com_byte_count(2), QN => spi_com_n_2);
  spi_com_byte_count_reg_3 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN322_spi_com_n_257, Q => spi_com_byte_count(3), QN => spi_com_n_4);
  spi_com_pause_count_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN279_spi_com_n_256, Q => spi_com_pause_count(2), QN => spi_com_n_8);
  spi_com_state_reg_0 : DFD1BWP7T port map(CP => CTS_19, D => spi_com_n_263, Q => spi_com_state(0), QN => spi_com_n_3);
  spi_com_drc_bufs11291 : INVD5BWP7T port map(I => spi_com_n_1, ZN => MOSI);
  spi_com_g2 : INR3D0BWP7T port map(A1 => spi_com_n_132, B1 => spi_com_n_19, B2 => spi_com_bit_count(2), ZN => spi_com_n_0);
  spi_com_state_reg_1 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN351_spi_com_n_254, Q => spi_com_state(1), QN => spi_com_n_264);
  spi_com_send_in0_reg : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => send, Q => spi_com_send_in0, QN => spi_com_n_10);

end routed;
