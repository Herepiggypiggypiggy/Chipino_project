
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of not_arduino is

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR4XD1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OA32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AO33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OA33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKSND1BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component CKAN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKND0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OA21D1BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  signal MISO_shift : std_logic_vector(72 downto 0);
  signal MOSI_shift : std_logic_vector(16 downto 0);
  signal full_map_2_2 : std_logic_vector(2 downto 0);
  signal full_map_9_14 : std_logic_vector(2 downto 0);
  signal full_map_5_2 : std_logic_vector(2 downto 0);
  signal full_map_2_0 : std_logic_vector(2 downto 0);
  signal full_map_2_14 : std_logic_vector(2 downto 0);
  signal full_map_1_13 : std_logic_vector(2 downto 0);
  signal full_map_2_1 : std_logic_vector(2 downto 0);
  signal full_map_0_14 : std_logic_vector(2 downto 0);
  signal full_map_10_11 : std_logic_vector(2 downto 0);
  signal full_map_0_13 : std_logic_vector(2 downto 0);
  signal full_map_3_2 : std_logic_vector(2 downto 0);
  signal full_map_3_5 : std_logic_vector(2 downto 0);
  signal full_map_4_0 : std_logic_vector(2 downto 0);
  signal full_map_14_13 : std_logic_vector(2 downto 0);
  signal full_map_14_11 : std_logic_vector(2 downto 0);
  signal full_map_14_1 : std_logic_vector(2 downto 0);
  signal full_map_4_1 : std_logic_vector(2 downto 0);
  signal full_map_6_2 : std_logic_vector(2 downto 0);
  signal full_map_1_2 : std_logic_vector(2 downto 0);
  signal full_map_0_5 : std_logic_vector(2 downto 0);
  signal full_map_6_0 : std_logic_vector(2 downto 0);
  signal full_map_5_14 : std_logic_vector(2 downto 0);
  signal full_map_0_2 : std_logic_vector(2 downto 0);
  signal full_map_1_1 : std_logic_vector(2 downto 0);
  signal full_map_14_12 : std_logic_vector(2 downto 0);
  signal full_map_4_2 : std_logic_vector(2 downto 0);
  signal full_map_14_14 : std_logic_vector(2 downto 0);
  signal full_map_14_2 : std_logic_vector(2 downto 0);
  signal full_map_1_0 : std_logic_vector(2 downto 0);
  signal full_map_0_4 : std_logic_vector(2 downto 0);
  signal full_map_12_14 : std_logic_vector(2 downto 0);
  signal full_map_5_0 : std_logic_vector(2 downto 0);
  signal full_map_3_14 : std_logic_vector(2 downto 0);
  signal full_map_4_14 : std_logic_vector(2 downto 0);
  signal full_map_0_12 : std_logic_vector(2 downto 0);
  signal full_map_1_14 : std_logic_vector(2 downto 0);
  signal full_map_0_11 : std_logic_vector(2 downto 0);
  signal full_map_6_14 : std_logic_vector(2 downto 0);
  signal full_map_3_0 : std_logic_vector(2 downto 0);
  signal full_map_0_9 : std_logic_vector(2 downto 0);
  signal full_map_14_10 : std_logic_vector(2 downto 0);
  signal full_map_0_3 : std_logic_vector(2 downto 0);
  signal full_map_8_12 : std_logic_vector(2 downto 0);
  signal full_map_0_1 : std_logic_vector(2 downto 0);
  signal full_map_0_0 : std_logic_vector(2 downto 0);
  signal full_map_14_0 : std_logic_vector(2 downto 0);
  signal full_map_14_4 : std_logic_vector(2 downto 0);
  signal full_map_14_3 : std_logic_vector(2 downto 0);
  signal full_map_10_14 : std_logic_vector(2 downto 0);
  signal full_map_9_0 : std_logic_vector(2 downto 0);
  signal full_map_7_10 : std_logic_vector(2 downto 0);
  signal full_map_11_4 : std_logic_vector(2 downto 0);
  signal full_map_14_5 : std_logic_vector(2 downto 0);
  signal full_map_11_0 : std_logic_vector(2 downto 0);
  signal full_map_13_0 : std_logic_vector(2 downto 0);
  signal full_map_7_0 : std_logic_vector(2 downto 0);
  signal full_map_8_0 : std_logic_vector(2 downto 0);
  signal full_map_5_6 : std_logic_vector(2 downto 0);
  signal full_map_0_10 : std_logic_vector(2 downto 0);
  signal full_map_0_6 : std_logic_vector(2 downto 0);
  signal full_map_0_8 : std_logic_vector(2 downto 0);
  signal full_map_0_7 : std_logic_vector(2 downto 0);
  signal full_map_12_0 : std_logic_vector(2 downto 0);
  signal full_map_8_4 : std_logic_vector(2 downto 0);
  signal full_map_10_0 : std_logic_vector(2 downto 0);
  signal full_map_14_6 : std_logic_vector(2 downto 0);
  signal full_map_11_14 : std_logic_vector(2 downto 0);
  signal full_map_8_14 : std_logic_vector(2 downto 0);
  signal full_map_14_9 : std_logic_vector(2 downto 0);
  signal full_map_10_8 : std_logic_vector(2 downto 0);
  signal full_map_10_12 : std_logic_vector(2 downto 0);
  signal full_map_7_14 : std_logic_vector(2 downto 0);
  signal full_map_13_14 : std_logic_vector(2 downto 0);
  signal full_map_14_8 : std_logic_vector(2 downto 0);
  signal full_map_14_7 : std_logic_vector(2 downto 0);
  signal bit_counter : std_logic_vector(3 downto 0);
  signal state : std_logic_vector(1 downto 0);
  signal UNCONNECTED, n_0, n_1, n_2, n_3 : std_logic;
  signal n_4, n_5, n_6, n_7, n_8 : std_logic;
  signal n_9, n_10, n_11, n_12, n_13 : std_logic;
  signal n_14, n_15, n_16, n_17, n_18 : std_logic;
  signal n_20, n_21, n_22, n_23, n_24 : std_logic;
  signal n_25, n_26, n_27, n_28, n_29 : std_logic;
  signal n_30, n_31, n_32, n_34, n_35 : std_logic;
  signal n_36, n_37, n_38, n_39, n_40 : std_logic;
  signal n_41, n_42, n_43, n_44, n_45 : std_logic;
  signal n_46, n_47, n_48, n_49, n_50 : std_logic;
  signal n_51, n_52, n_53, n_54, n_55 : std_logic;
  signal n_56, n_57, n_58, n_59, n_60 : std_logic;
  signal n_61, n_62, n_63, n_64, n_65 : std_logic;
  signal n_66, n_67, n_68, n_69, n_70 : std_logic;
  signal n_71, n_72, n_73, n_74, n_75 : std_logic;
  signal n_76, n_77, n_78, n_79, n_80 : std_logic;
  signal n_81, n_82, n_83, n_84, n_85 : std_logic;
  signal n_86, n_87, n_88, n_89, n_90 : std_logic;
  signal n_91, n_92, n_93, n_94, n_95 : std_logic;
  signal n_96, n_97, n_98, n_99, n_100 : std_logic;
  signal n_101, n_102, n_103, n_104, n_105 : std_logic;
  signal n_106, n_107, n_108, n_109, n_110 : std_logic;
  signal n_111, n_112, n_113, n_114, n_115 : std_logic;
  signal n_116, n_117, n_118, n_119, n_121 : std_logic;
  signal n_122, n_123, n_124, n_125, n_126 : std_logic;
  signal n_127, n_128, n_129, n_130, n_131 : std_logic;
  signal n_132, n_133, n_134, n_135, n_136 : std_logic;
  signal n_137, n_138, n_139, n_140, n_141 : std_logic;
  signal n_142, n_143, n_144, n_145, n_146 : std_logic;
  signal n_147, n_148, n_149, n_150, n_151 : std_logic;
  signal n_152, n_153, n_154, n_155, n_156 : std_logic;
  signal n_157, n_158, n_159, n_160, n_161 : std_logic;
  signal n_162, n_164, n_165, n_166, n_167 : std_logic;
  signal n_168, n_169, n_170, n_171, n_172 : std_logic;
  signal n_173, n_174, n_175, n_176, n_177 : std_logic;
  signal n_178, n_179, n_180, n_181, n_182 : std_logic;
  signal n_183, n_184, n_185, n_186, n_187 : std_logic;
  signal n_188, n_189, n_190, n_191, n_192 : std_logic;
  signal n_193, n_194, n_195, n_196, n_197 : std_logic;
  signal n_198, n_199, n_200, n_201, n_202 : std_logic;
  signal n_203, n_204, n_205, n_206, n_207 : std_logic;
  signal n_208, n_209, n_210, n_211, n_212 : std_logic;
  signal n_213, n_214, n_215, n_216, n_217 : std_logic;
  signal n_218, n_219, n_220, n_221, n_222 : std_logic;
  signal n_223, n_224, n_225, n_226, n_227 : std_logic;
  signal n_228, n_229, n_230, n_231, n_232 : std_logic;
  signal n_233, n_234, n_235, n_236, n_237 : std_logic;
  signal n_238, n_239, n_240, n_241, n_242 : std_logic;
  signal n_243, n_244, n_245, n_246, n_247 : std_logic;
  signal n_248, n_249, n_250, n_251, n_252 : std_logic;
  signal n_253, n_254, n_255, n_256, n_257 : std_logic;
  signal n_258, n_259, n_260, n_261, n_262 : std_logic;
  signal n_263, n_264, n_265, n_266, n_267 : std_logic;
  signal n_268, n_269, n_270, n_271, n_272 : std_logic;
  signal n_273, n_274, n_275, n_276, n_277 : std_logic;
  signal n_278, n_279, n_280, n_281, n_282 : std_logic;
  signal n_283, n_284, n_285, n_286, n_287 : std_logic;
  signal n_288, n_289, n_290, n_291, n_292 : std_logic;
  signal n_293, n_294, n_295, n_296, n_297 : std_logic;
  signal n_298, n_299, n_300, n_301, n_302 : std_logic;
  signal n_303, n_304, n_305, n_306, n_307 : std_logic;
  signal n_308, n_309, n_310, n_311, n_312 : std_logic;
  signal n_313, n_314, n_315, n_316, n_317 : std_logic;
  signal n_318, n_319, n_320, n_321, n_322 : std_logic;
  signal n_323, n_324, n_325, n_326, n_327 : std_logic;
  signal n_328, n_329, n_330, n_332, n_333 : std_logic;
  signal n_334, n_335, n_336, n_337, n_338 : std_logic;
  signal n_339, n_340, n_341, n_342, n_343 : std_logic;
  signal n_344, n_345, n_346, n_347, n_348 : std_logic;
  signal n_349, n_350, n_351, n_352, n_353 : std_logic;
  signal n_354, n_355, n_356, n_357, n_358 : std_logic;
  signal n_359, n_360, n_361, n_362, n_363 : std_logic;
  signal n_364, n_365, n_366, n_367, n_368 : std_logic;
  signal n_369, n_370, n_371, n_372, n_373 : std_logic;
  signal n_374, n_375, n_376, n_377, n_379 : std_logic;
  signal n_380, n_381, n_382, n_383, n_384 : std_logic;
  signal n_385, n_386, n_387, n_388, n_389 : std_logic;
  signal n_390, n_391, n_392, n_393, n_394 : std_logic;
  signal n_395, n_396, n_397, n_398, n_399 : std_logic;
  signal n_400, n_401, n_402, n_403, n_404 : std_logic;
  signal n_405, n_406, n_407, n_408, n_409 : std_logic;
  signal n_410, n_411, n_412, n_413, n_414 : std_logic;
  signal n_415, n_416, n_417, n_418, n_419 : std_logic;
  signal n_420, n_421, n_422, n_423, n_424 : std_logic;
  signal n_425, n_426, n_427, n_428, n_429 : std_logic;
  signal n_430, n_431, n_432, n_433, n_434 : std_logic;
  signal n_435, n_436, n_437, n_438, n_439 : std_logic;
  signal n_440, n_441, n_442, n_443, n_444 : std_logic;
  signal n_445, n_446, n_447, n_448, n_449 : std_logic;
  signal n_450, n_451, n_452, n_453, n_454 : std_logic;
  signal n_455, n_456, n_457, n_458, n_459 : std_logic;
  signal n_460, n_461, n_462, n_463, n_464 : std_logic;
  signal n_465, n_466, n_467, n_468, n_469 : std_logic;
  signal n_470, n_471, n_472, n_473, n_474 : std_logic;
  signal n_475, n_476, n_477, n_478, n_479 : std_logic;
  signal n_480, n_481, n_482, n_483, n_484 : std_logic;
  signal n_485, n_486, n_487, n_488, n_489 : std_logic;
  signal n_490, n_491, n_492, n_493, n_494 : std_logic;
  signal n_495, n_496, n_497, n_498, n_499 : std_logic;
  signal n_500, n_501, n_502, n_503, n_504 : std_logic;
  signal n_505, n_506, n_507, n_508, n_509 : std_logic;
  signal n_510, n_511, n_512, n_513, n_514 : std_logic;
  signal n_515, n_516, n_517, n_518, n_519 : std_logic;
  signal n_520, n_521, n_522, n_523, n_524 : std_logic;
  signal n_525, n_526, n_527, n_528, n_529 : std_logic;
  signal n_530, n_531, n_532, n_533, n_534 : std_logic;
  signal n_535, n_536, n_537, n_538, n_539 : std_logic;
  signal n_540, n_541, n_542, n_543, n_544 : std_logic;
  signal n_545, n_546, n_547, n_548, n_549 : std_logic;
  signal n_550, n_551, n_552, n_553, n_554 : std_logic;
  signal n_555, n_556, n_557, n_558, n_559 : std_logic;
  signal n_560, n_561, n_562, n_563, n_564 : std_logic;
  signal n_565, n_566, n_567, n_568, n_569 : std_logic;
  signal n_570, n_571, n_572, n_573, n_574 : std_logic;
  signal n_575, n_576, n_577, n_578, n_579 : std_logic;
  signal n_580, n_581, n_582, n_583, n_584 : std_logic;
  signal n_585, n_586, n_587, n_588, n_589 : std_logic;
  signal n_590, n_591, n_592, n_593, n_594 : std_logic;
  signal n_595, n_596, n_597, n_598, n_599 : std_logic;
  signal n_600, n_601, n_602, n_603, n_604 : std_logic;
  signal n_605, n_606, n_607, n_608, n_609 : std_logic;
  signal n_610, n_611, n_612, n_613, n_614 : std_logic;
  signal n_615, n_616, n_617, n_618, n_619 : std_logic;
  signal n_620, n_621, n_622, n_623, n_624 : std_logic;
  signal n_625, n_626, n_627, n_628, n_629 : std_logic;
  signal n_630, n_631, n_632, n_633, n_634 : std_logic;
  signal n_635, n_636, n_637, n_638, n_639 : std_logic;
  signal n_640, n_641, n_642, n_643, n_644 : std_logic;
  signal n_645, n_646, n_647, n_648, n_649 : std_logic;
  signal n_650, n_651, n_652, n_653, n_654 : std_logic;
  signal n_655, n_656, n_657, n_658, n_659 : std_logic;
  signal n_660, n_661, n_662, n_663, n_664 : std_logic;
  signal n_665, n_666, n_667, n_668, n_669 : std_logic;
  signal n_670, n_671, n_672, n_673, n_674 : std_logic;
  signal n_675, n_676, n_677, n_678, n_679 : std_logic;
  signal n_680, n_681, n_682, n_683, n_684 : std_logic;
  signal n_685, n_686, n_687, n_688, n_689 : std_logic;
  signal n_690, n_691, n_692, n_693, n_694 : std_logic;
  signal n_695, n_696, n_697, n_698, n_699 : std_logic;
  signal n_700, n_701, n_702, n_703, n_704 : std_logic;
  signal n_705, n_706, n_707, n_708, n_709 : std_logic;
  signal n_710, n_711, n_712, n_713, n_714 : std_logic;
  signal n_715, n_716, n_717, n_718, n_719 : std_logic;
  signal n_720, n_721, n_722, n_723, n_724 : std_logic;
  signal n_725, n_726, n_727, n_728, n_729 : std_logic;
  signal n_730, n_731, n_732, n_733, n_734 : std_logic;
  signal n_735, n_736, n_737, n_738, n_739 : std_logic;
  signal n_740, n_741, n_742, n_743, n_744 : std_logic;
  signal n_745, n_746, n_747, n_748, n_749 : std_logic;
  signal n_750, n_751, n_752, n_753, n_754 : std_logic;
  signal n_755, n_756, n_757, n_758, n_759 : std_logic;
  signal n_760, n_761, n_762, n_763, n_764 : std_logic;
  signal n_765, n_766, n_767, n_768, n_769 : std_logic;
  signal n_770, n_771, n_772, n_773, n_774 : std_logic;
  signal n_775, n_776, n_777, n_778, n_779 : std_logic;
  signal n_780, n_781, n_782, n_783, n_784 : std_logic;
  signal n_785, n_786, n_787, n_788, n_789 : std_logic;
  signal n_790, n_791, n_792, n_793, n_794 : std_logic;
  signal n_795, n_796, n_797, n_798, n_799 : std_logic;
  signal n_800, n_801, n_802, n_803, n_804 : std_logic;
  signal n_805, n_806, n_807, n_808, n_809 : std_logic;
  signal n_810, n_811, n_812, n_813, n_814 : std_logic;
  signal n_815, n_816, n_817, n_818, n_819 : std_logic;
  signal n_820, n_821, n_822, n_823, n_824 : std_logic;
  signal n_825, n_826, n_827, n_828, n_829 : std_logic;
  signal n_830, n_831, n_832, n_833, n_834 : std_logic;
  signal n_835, n_836, n_837, n_838, n_839 : std_logic;
  signal n_840, n_841, n_842, n_843, n_844 : std_logic;
  signal n_845, n_846, n_847, n_848, n_849 : std_logic;
  signal n_850, n_851, n_852, n_853, n_854 : std_logic;
  signal n_855, n_856, n_857, n_858, n_859 : std_logic;
  signal n_860, n_861, n_862, n_863, n_864 : std_logic;
  signal n_865, n_866, n_867, n_868, n_869 : std_logic;
  signal n_870, n_871, n_872, n_873, n_874 : std_logic;
  signal n_875, n_876, n_877, n_878, n_879 : std_logic;
  signal n_880, n_881, n_882, n_883, n_884 : std_logic;
  signal n_885, n_886, n_887, n_888, n_889 : std_logic;
  signal n_890, n_891, n_892, n_893, n_894 : std_logic;
  signal n_895, n_896, n_897, n_898, n_899 : std_logic;
  signal n_900, n_901, n_902, n_903, n_904 : std_logic;
  signal n_905, n_906, n_907, n_908, n_909 : std_logic;
  signal n_910, n_911, n_912, n_913, n_914 : std_logic;
  signal n_915, n_916, n_917, n_918, n_919 : std_logic;
  signal n_920, n_921, n_922, n_923, n_924 : std_logic;
  signal n_925, n_926, n_927, n_928, n_929 : std_logic;
  signal n_930, n_932, n_933, n_934, n_935 : std_logic;
  signal n_936, n_937, n_938, n_939, n_940 : std_logic;
  signal n_941, n_942, n_943, n_944, n_945 : std_logic;
  signal n_946, n_947, n_948, n_949, n_950 : std_logic;
  signal n_951, n_952, n_953, n_954, n_955 : std_logic;
  signal n_956, n_957, n_958, n_959, n_960 : std_logic;
  signal n_961, n_962, n_963, n_964, n_965 : std_logic;
  signal n_966, n_967, n_968, n_969, n_970 : std_logic;
  signal n_971, n_972, n_973, n_974, n_975 : std_logic;
  signal n_976, n_977, n_978, n_979, n_980 : std_logic;
  signal n_981, n_982, n_983, n_985, n_986 : std_logic;
  signal n_987, n_988, n_989, n_990, n_991 : std_logic;
  signal n_992, n_993, n_994, n_995, n_996 : std_logic;
  signal n_997, n_998, n_999, n_1000, n_1001 : std_logic;
  signal n_1002, n_1003, n_1004, n_1005, n_1006 : std_logic;
  signal n_1007, n_1008, n_1009, n_1010, n_1011 : std_logic;
  signal n_1012, n_1013, n_1014, n_1015, n_1016 : std_logic;
  signal n_1017, n_1018, n_1019, n_1020, n_1021 : std_logic;
  signal n_1022, n_1023, n_1024, n_1025, n_1026 : std_logic;
  signal n_1027, n_1028, n_1029, n_1030, n_1031 : std_logic;
  signal n_1032, n_1033, n_1034, n_1035, n_1036 : std_logic;
  signal n_1037, n_1038, n_1039, n_1040, n_1041 : std_logic;
  signal n_1042, n_1043, n_1044, n_1045, n_1046 : std_logic;
  signal n_1047, n_1048, n_1049, n_1050, n_1052 : std_logic;
  signal n_1053, n_1054, n_1055, n_1056, n_1057 : std_logic;
  signal n_1058, n_1059, n_1060, n_1061, n_1062 : std_logic;
  signal n_1063, n_1064, n_1065, n_1066, n_1067 : std_logic;
  signal n_1068, n_1069, n_1070, n_1071, n_1072 : std_logic;
  signal n_1073, n_1074, n_1075, n_1076, n_1077 : std_logic;
  signal n_1078, n_1079, n_1080, n_1081, n_1082 : std_logic;
  signal n_1083, n_1084, n_1085, n_1086, n_1087 : std_logic;
  signal n_1088, n_1089, n_1090, n_1091, n_1092 : std_logic;
  signal n_1093, n_1094, n_1095, n_1096, n_1097 : std_logic;
  signal n_1098, n_1099, n_1100, n_1101, n_1102 : std_logic;
  signal n_1103, n_1104, n_1105, n_1106, n_1107 : std_logic;
  signal n_1108, n_1109, n_1110, n_1111, n_1112 : std_logic;
  signal n_1113, n_1114, n_1115, n_1116, n_1117 : std_logic;
  signal n_1118, n_1119, n_1120, n_1121, n_1122 : std_logic;
  signal n_1123, n_1124, n_1125, n_1126, n_1127 : std_logic;
  signal n_1128, n_1129, n_1130, n_1131, n_1132 : std_logic;
  signal n_1133, n_1134, n_1135, n_1136, n_1137 : std_logic;
  signal n_1138, n_1139, n_1140, n_1141, n_1142 : std_logic;
  signal n_1143, n_1144, n_1145, n_1146, n_1147 : std_logic;
  signal n_1148, n_1149, n_1150, n_1151, n_1152 : std_logic;
  signal n_1153, n_1154, n_1155, n_1156, n_1157 : std_logic;
  signal n_1158, n_1159, n_1160, n_1161, n_1162 : std_logic;
  signal n_1163, n_1164, n_1165, n_1166, n_1167 : std_logic;
  signal n_1168, n_1169, n_1170, n_1171, n_1172 : std_logic;
  signal n_1173, n_1174, n_1175, n_1176, n_1177 : std_logic;
  signal n_1178, n_1179, n_1180, n_1181, n_1182 : std_logic;
  signal n_1183, n_1184, n_1185, n_1187, n_1188 : std_logic;
  signal n_1189, n_1190, n_1191, n_1192, n_1193 : std_logic;
  signal n_1194, n_1195, n_1196, n_1197, n_1198 : std_logic;
  signal n_1199, n_1200, n_1201, n_1202, n_1203 : std_logic;
  signal n_1204, n_1205, n_1206, n_1207, n_1208 : std_logic;
  signal n_1209, n_1210, n_1211, n_1212, n_1213 : std_logic;
  signal n_1214, n_1215, n_1216, n_1217, n_1218 : std_logic;
  signal n_1219, n_1220, n_1221, n_1222, n_1223 : std_logic;
  signal n_1224, n_1225, n_1226, n_1227, n_1228 : std_logic;
  signal n_1229, n_1230, n_1231, n_1232, n_1233 : std_logic;
  signal n_1234, n_1235, n_1236, n_1237, n_1238 : std_logic;
  signal n_1239, n_1240, n_1241, n_1242, n_1243 : std_logic;
  signal n_1244, n_1252, n_1256, n_1257, n_1258 : std_logic;
  signal n_1259, n_1260 : std_logic;

begin

  MISO_shift_reg_10 : DFQD1BWP7T port map(CP => clk, D => n_1243, Q => MISO_shift(10));
  MISO_shift_reg_70 : DFQD1BWP7T port map(CP => clk, D => n_1241, Q => MISO_shift(70));
  MISO_shift_reg_55 : DFQD1BWP7T port map(CP => clk, D => n_1244, Q => MISO_shift(55));
  MISO_shift_reg_46 : DFQD1BWP7T port map(CP => clk, D => n_1240, Q => MISO_shift(46));
  MISO_shift_reg_34 : DFQD1BWP7T port map(CP => clk, D => n_1238, Q => MISO_shift(34));
  MISO_shift_reg_13 : DFQD1BWP7T port map(CP => clk, D => n_1237, Q => MISO_shift(13));
  g89068 : ND4D0BWP7T port map(A1 => n_1222, A2 => n_1217, A3 => n_1239, A4 => n_1242, ZN => n_1244);
  g89059 : ND4D0BWP7T port map(A1 => n_1228, A2 => n_1115, A3 => n_1231, A4 => n_1242, ZN => n_1243);
  MISO_shift_reg_28 : DFQD1BWP7T port map(CP => clk, D => n_1235, Q => MISO_shift(28));
  g89060 : ND4D0BWP7T port map(A1 => n_1227, A2 => n_975, A3 => n_974, A4 => n_1224, ZN => n_1241);
  MISO_shift_reg_4 : DFQD1BWP7T port map(CP => clk, D => n_1233, Q => MISO_shift(4));
  MISO_shift_reg_52 : DFQD1BWP7T port map(CP => clk, D => n_1230, Q => MISO_shift(52));
  MISO_shift_reg_19 : DFQD1BWP7T port map(CP => clk, D => n_1234, Q => MISO_shift(19));
  g89057 : ND3D0BWP7T port map(A1 => n_1223, A2 => n_1239, A3 => n_1236, ZN => n_1240);
  g89051 : IND4D0BWP7T port map(A1 => n_1135, B1 => n_1232, B2 => n_1192, B3 => n_1213, ZN => n_1238);
  g89069 : ND2D1BWP7T port map(A1 => n_1226, A2 => n_1236, ZN => n_1237);
  MISO_shift_reg_67 : DFQD1BWP7T port map(CP => clk, D => n_1225, Q => MISO_shift(67));
  MISO_shift_reg_31 : DFQD1BWP7T port map(CP => clk, D => n_1221, Q => MISO_shift(31));
  MISO_shift_reg_37 : DFQD1BWP7T port map(CP => clk, D => n_1229, Q => MISO_shift(37));
  g89056 : ND3D0BWP7T port map(A1 => n_1219, A2 => n_1144, A3 => n_1143, ZN => n_1235);
  g89105 : IND4D0BWP7T port map(A1 => n_970, B1 => n_1215, B2 => n_1084, B3 => n_1211, ZN => n_1234);
  g89082 : IND4D0BWP7T port map(A1 => n_1206, B1 => n_1232, B2 => n_1231, B3 => n_1043, ZN => n_1233);
  g89087 : ND3D0BWP7T port map(A1 => n_1220, A2 => n_1181, A3 => n_1239, ZN => n_1230);
  MISO_shift_reg_22 : DFQD1BWP7T port map(CP => clk, D => n_1216, Q => MISO_shift(22));
  MISO_shift_reg_17 : DFQD1BWP7T port map(CP => clk, D => n_1214, Q => MISO_shift(17));
  MISO_shift_reg_56 : DFQD1BWP7T port map(CP => clk, D => n_1218, Q => MISO_shift(56));
  g89104 : IND4D0BWP7T port map(A1 => n_1066, B1 => n_1242, B2 => n_1160, B3 => n_1201, ZN => n_1229);
  g89101 : NR4D0BWP7T port map(A1 => n_1199, A2 => n_983, A3 => n_1113, A4 => n_1114, ZN => n_1228);
  g89100 : NR4D0BWP7T port map(A1 => n_1202, A2 => n_891, A3 => n_890, A4 => n_889, ZN => n_1227);
  g89083 : NR4D0BWP7T port map(A1 => n_1189, A2 => n_1111, A3 => n_1110, A4 => n_1109, ZN => n_1226);
  g89067 : ND4D0BWP7T port map(A1 => n_1205, A2 => n_1033, A3 => n_1224, A4 => n_1242, ZN => n_1225);
  g89085 : NR4D0BWP7T port map(A1 => n_1197, A2 => n_1122, A3 => n_1121, A4 => n_1190, ZN => n_1223);
  g89120 : INR4D0BWP7T port map(A1 => n_1125, B1 => n_1177, B2 => n_1178, B3 => n_1196, ZN => n_1222);
  g89073 : ND2D0BWP7T port map(A1 => n_1212, A2 => n_1236, ZN => n_1221);
  MISO_shift_reg_32 : DFQD1BWP7T port map(CP => clk, D => n_1210, Q => MISO_shift(32));
  MISO_shift_reg_16 : DFQD1BWP7T port map(CP => clk, D => n_1209, Q => MISO_shift(16));
  MISO_shift_reg_25 : DFQD1BWP7T port map(CP => clk, D => n_1207, Q => MISO_shift(25));
  g89122 : NR4D0BWP7T port map(A1 => n_1180, A2 => n_1182, A3 => n_1100, A4 => n_1099, ZN => n_1220);
  g89086 : NR4D0BWP7T port map(A1 => n_1187, A2 => n_1037, A3 => n_1036, A4 => n_1035, ZN => n_1219);
  g89119 : ND4D0BWP7T port map(A1 => n_1179, A2 => n_1217, A3 => n_1239, A4 => n_1242, ZN => n_1218);
  g89088 : IND4D0BWP7T port map(A1 => n_1173, B1 => n_1242, B2 => n_1215, B3 => n_1140, ZN => n_1216);
  g89125 : ND4D0BWP7T port map(A1 => n_1188, A2 => n_1208, A3 => n_1215, A4 => n_1232, ZN => n_1214);
  g89093 : NR3D0BWP7T port map(A1 => n_1198, A2 => n_1193, A3 => n_732, ZN => n_1213);
  MISO_shift_reg_49 : DFQD1BWP7T port map(CP => clk, D => n_1195, Q => MISO_shift(49));
  MISO_shift_reg_23 : DFQD1BWP7T port map(CP => clk, D => n_1200, Q => MISO_shift(23));
  MISO_shift_reg_58 : DFQD1BWP7T port map(CP => clk, D => n_1204, Q => MISO_shift(58));
  MISO_shift_reg_35 : DFQD1BWP7T port map(CP => clk, D => n_1194, Q => MISO_shift(35));
  MISO_shift_reg_47 : DFQD1BWP7T port map(CP => clk, D => n_1191, Q => MISO_shift(47));
  g89102 : NR4D0BWP7T port map(A1 => n_1166, A2 => n_1171, A3 => n_1170, A4 => n_1169, ZN => n_1212);
  g89155 : INR4D0BWP7T port map(A1 => n_1083, B1 => n_918, B2 => n_969, B3 => n_1158, ZN => n_1211);
  g89118 : ND2D0BWP7T port map(A1 => n_1172, A2 => n_1236, ZN => n_1210);
  g89090 : ND4D0BWP7T port map(A1 => n_1156, A2 => n_1208, A3 => n_1215, A4 => n_1232, ZN => n_1209);
  MISO_shift_reg_14 : DFQD1BWP7T port map(CP => clk, D => n_1185, Q => MISO_shift(14));
  MISO_shift_reg_1 : DFQD1BWP7T port map(CP => clk, D => n_1176, Q => MISO_shift(1));
  g89071 : IND4D0BWP7T port map(A1 => n_937, B1 => n_1203, B2 => n_1054, B3 => n_1162, ZN => n_1207);
  g89142 : ND4D0BWP7T port map(A1 => n_1157, A2 => n_1127, A3 => n_850, A4 => n_1042, ZN => n_1206);
  MISO_shift_reg_7 : DFQD1BWP7T port map(CP => clk, D => n_1174, Q => MISO_shift(7));
  MISO_shift_reg_53 : DFQD1BWP7T port map(CP => clk, D => n_1183, Q => MISO_shift(53));
  MISO_shift_reg_11 : DFQD1BWP7T port map(CP => clk, D => n_1256, Q => MISO_shift(11));
  MISO_shift_reg_43 : DFQD1BWP7T port map(CP => clk, D => n_1175, Q => MISO_shift(43));
  g89109 : NR3D0BWP7T port map(A1 => n_1167, A2 => n_1031, A3 => n_1032, ZN => n_1205);
  g89106 : IND4D0BWP7T port map(A1 => n_1137, B1 => n_1203, B2 => n_1239, B3 => n_1102, ZN => n_1204);
  g89158 : IND4D0BWP7T port map(A1 => n_608, B1 => n_617, B2 => n_607, B3 => n_1151, ZN => n_1202);
  g89160 : AN4D0BWP7T port map(A1 => n_1148, A2 => n_963, A3 => n_885, A4 => n_1159, Z => n_1201);
  g89108 : ND4D0BWP7T port map(A1 => n_1141, A2 => n_1096, A3 => n_1215, A4 => n_1242, ZN => n_1200);
  g89162 : OAI211D1BWP7T port map(A1 => n_1117, A2 => n_995, B => n_1120, C => n_685, ZN => n_1199);
  g89149 : AO221D0BWP7T port map(A1 => n_962, A2 => n_1015, B1 => n_1089, B2 => n_1092, C => n_1165, Z => n_1198);
  g89131 : IND3D0BWP7T port map(A1 => n_1029, B1 => n_1123, B2 => n_1134, ZN => n_1197);
  g89182 : ND4D0BWP7T port map(A1 => n_1149, A2 => n_879, A3 => n_740, A4 => n_719, ZN => n_1196);
  g89089 : IND4D0BWP7T port map(A1 => n_1072, B1 => n_1232, B2 => n_1239, B3 => n_1130, ZN => n_1195);
  g89126 : IND4D0BWP7T port map(A1 => n_1193, B1 => n_1232, B2 => n_1192, B3 => n_1136, ZN => n_1194);
  g89084 : IND4D0BWP7T port map(A1 => n_1190, B1 => n_1236, B2 => n_1239, B3 => n_1124, ZN => n_1191);
  g89132 : ND3D0BWP7T port map(A1 => n_1164, A2 => n_1000, A3 => n_1184, ZN => n_1189);
  MISO_shift_reg_38 : DFQD1BWP7T port map(CP => clk, D => n_1161, Q => MISO_shift(38));
  MISO_shift_reg_50 : DFQD1BWP7T port map(CP => clk, D => n_1168, Q => MISO_shift(50));
  g89167 : NR4D0BWP7T port map(A1 => n_1118, A2 => n_1155, A3 => n_1154, A4 => n_1153, ZN => n_1188);
  g89147 : ND4D0BWP7T port map(A1 => n_1104, A2 => n_949, A3 => n_615, A4 => n_1142, ZN => n_1187);
  g89107 : ND4D0BWP7T port map(A1 => n_1112, A2 => n_1184, A3 => n_1163, A4 => n_1236, ZN => n_1185);
  g89144 : IND4D0BWP7T port map(A1 => n_1182, B1 => n_1239, B2 => n_1181, B3 => n_1101, ZN => n_1183);
  g89168 : IND4D0BWP7T port map(A1 => n_1106, B1 => n_757, B2 => n_840, B3 => n_914, ZN => n_1180);
  g89170 : NR3D0BWP7T port map(A1 => n_1126, A2 => n_1178, A3 => n_1177, ZN => n_1179);
  g89058 : ND2D1BWP7T port map(A1 => n_1133, A2 => n_1231, ZN => n_1176);
  g89092 : IND4D0BWP7T port map(A1 => n_1119, B1 => n_1063, B2 => n_922, B3 => n_923, ZN => n_1175);
  g89091 : IND4D0BWP7T port map(A1 => n_1047, B1 => n_1231, B2 => n_1094, B3 => n_1098, ZN => n_1174);
  g89130 : IND4D0BWP7T port map(A1 => n_1139, B1 => n_1039, B2 => n_1040, B3 => n_1097, ZN => n_1173);
  g89140 : NR4D0BWP7T port map(A1 => n_1105, A2 => n_1171, A3 => n_1170, A4 => n_1169, ZN => n_1172);
  MISO_shift_reg_64 : DFQD1BWP7T port map(CP => clk, D => n_1152, Q => MISO_shift(64));
  MISO_shift_reg_5 : DFQD1BWP7T port map(CP => clk, D => n_1128, Q => MISO_shift(5));
  MISO_shift_reg_2 : DFQD1BWP7T port map(CP => clk, D => n_1138, Q => MISO_shift(2));
  MISO_shift_reg_29 : DFQD1BWP7T port map(CP => clk, D => n_1145, Q => MISO_shift(29));
  g89127 : ND4D0BWP7T port map(A1 => n_1075, A2 => n_1129, A3 => n_1239, A4 => n_1232, ZN => n_1168);
  g89159 : OAI211D1BWP7T port map(A1 => MOSI_shift(2), A2 => n_426, B => n_1061, C => n_397, ZN => n_1167);
  g89163 : ND4D0BWP7T port map(A1 => n_1088, A2 => n_930, A3 => n_900, A4 => n_374, ZN => n_1166);
  g89169 : OAI211D0BWP7T port map(A1 => n_1052, A2 => n_785, B => n_1082, C => n_561, ZN => n_1165);
  g89172 : INR3D0BWP7T port map(A1 => n_1163, B1 => n_1001, B2 => n_1071, ZN => n_1164);
  g89123 : NR4D0BWP7T port map(A1 => n_1078, A2 => n_939, A3 => n_938, A4 => n_1055, ZN => n_1162);
  g89146 : ND4D0BWP7T port map(A1 => n_1067, A2 => n_1160, A3 => n_1159, A4 => n_1242, ZN => n_1161);
  g89216 : ND4D0BWP7T port map(A1 => n_1093, A2 => n_934, A3 => n_689, A4 => n_473, ZN => n_1158);
  g89202 : AOI221D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(3), B1 => n_1091, B2 => n_1080, C => n_1079, ZN => n_1157);
  g89134 : NR4D0BWP7T port map(A1 => n_1069, A2 => n_1155, A3 => n_1154, A4 => n_1153, ZN => n_1156);
  MISO_shift_reg_59 : DFQD1BWP7T port map(CP => clk, D => n_1103, Q => MISO_shift(59));
  MISO_shift_reg_68 : DFQD1BWP7T port map(CP => clk, D => n_1107, Q => MISO_shift(68));
  MISO_shift_reg_40 : DFQD1BWP7T port map(CP => clk, D => n_1108, Q => MISO_shift(40));
  MISO_shift_reg_8 : DFQD1BWP7T port map(CP => clk, D => n_1095, Q => MISO_shift(8));
  g89143 : IND4D0BWP7T port map(A1 => n_1025, B1 => n_1224, B2 => n_1076, B3 => n_988, ZN => n_1152);
  g89221 : AOI221D0BWP7T port map(A1 => n_911, A2 => n_1086, B1 => n_1150, B2 => MISO_shift(69), C => n_1057, ZN => n_1151);
  g89224 : AOI22D0BWP7T port map(A1 => n_1147, A2 => n_1090, B1 => n_942, B2 => n_1146, ZN => n_1149);
  g89226 : AOI22D0BWP7T port map(A1 => n_1147, A2 => n_1146, B1 => n_878, B2 => n_1087, ZN => n_1148);
  g89148 : ND4D0BWP7T port map(A1 => n_1038, A2 => n_1144, A3 => n_1143, A4 => n_1142, ZN => n_1145);
  g89153 : INR3D0BWP7T port map(A1 => n_1140, B1 => n_1139, B2 => n_1041, ZN => n_1141);
  g89121 : OR4XD1BWP7T port map(A1 => n_869, A2 => n_1131, A3 => n_1132, A4 => n_1257, Z => n_1138);
  g89161 : ND3D0BWP7T port map(A1 => n_1070, A2 => n_998, A3 => n_997, ZN => n_1137);
  g89171 : NR3D0BWP7T port map(A1 => n_1060, A2 => n_882, A3 => n_1135, ZN => n_1136);
  MISO_shift_reg_44 : DFQD1BWP7T port map(CP => clk, D => n_1065, Q => MISO_shift(44));
  g89180 : NR4D0BWP7T port map(A1 => n_1058, A2 => n_783, A3 => n_695, A4 => n_1028, ZN => n_1134);
  g89070 : NR4D0BWP7T port map(A1 => n_1059, A2 => n_956, A3 => n_1132, A4 => n_1131, ZN => n_1133);
  g89129 : AN4D0BWP7T port map(A1 => n_1027, A2 => n_1129, A3 => n_1074, A4 => n_1073, Z => n_1130);
  g89141 : IND4D0BWP7T port map(A1 => n_1044, B1 => n_1232, B2 => n_1231, B3 => n_1127, ZN => n_1128);
  g89213 : ND4D0BWP7T port map(A1 => n_1049, A2 => n_868, A3 => n_1125, A4 => n_236, ZN => n_1126);
  g89139 : IINR4D0BWP7T port map(A1 => n_1030, A2 => n_1123, B1 => n_1122, B2 => n_1121, ZN => n_1124);
  g89207 : AOI211D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(9), B => n_1053, C => n_393, ZN => n_1120);
  MISO_shift_reg_65 : DFQD1BWP7T port map(CP => clk, D => n_1077, Q => MISO_shift(65));
  MISO_shift_reg_61 : DFQD1BWP7T port map(CP => clk, D => n_1068, Q => MISO_shift(61));
  MISO_shift_reg_20 : DFQD1BWP7T port map(CP => clk, D => n_1085, Q => MISO_shift(20));
  g89156 : IND3D0BWP7T port map(A1 => n_1064, B1 => n_1062, B2 => n_1005, ZN => n_1119);
  g89231 : OAI211D1BWP7T port map(A1 => n_1117, A2 => n_595, B => n_1023, C => n_503, ZN => n_1118);
  g89150 : INR4D0BWP7T port map(A1 => n_1115, B1 => n_1114, B2 => n_1113, B3 => n_1007, ZN => n_1116);
  g89151 : NR4D0BWP7T port map(A1 => n_1002, A2 => n_1111, A3 => n_1110, A4 => n_1109, ZN => n_1112);
  g89152 : IND3D0BWP7T port map(A1 => n_1003, B1 => n_1203, B2 => n_1006, ZN => n_1108);
  g89154 : ND3D0BWP7T port map(A1 => n_1034, A2 => n_1224, A3 => n_1242, ZN => n_1107);
  g89223 : OAI22D0BWP7T port map(A1 => n_1045, A2 => n_1010, B1 => n_724, B2 => n_781, ZN => n_1106);
  g89195 : OAI211D1BWP7T port map(A1 => n_965, A2 => n_883, B => n_1020, C => n_229, ZN => n_1105);
  g89205 : AOI211XD0BWP7T port map(A1 => n_1022, A2 => MISO_shift(28), B => n_1021, C => n_402, ZN => n_1104);
  g89166 : ND4D0BWP7T port map(A1 => n_999, A2 => n_1102, A3 => n_1239, A4 => n_1203, ZN => n_1103);
  g89184 : NR4D0BWP7T port map(A1 => n_951, A2 => n_1011, A3 => n_1100, A4 => n_1099, ZN => n_1101);
  g89164 : NR4D0BWP7T port map(A1 => n_996, A2 => n_835, A3 => n_1014, A4 => n_1046, ZN => n_1098);
  g89204 : AN4D0BWP7T port map(A1 => n_964, A2 => n_1008, A3 => n_821, A4 => n_1096, Z => n_1097);
  g89133 : ND3D0BWP7T port map(A1 => n_1048, A2 => n_1094, A3 => n_1231, ZN => n_1095);
  MISO_shift_reg_26 : DFQD1BWP7T port map(CP => clk, D => n_1056, Q => MISO_shift(26));
  g89274 : AOI222D0BWP7T port map(A1 => n_936, A2 => n_1092, B1 => n_1091, B2 => n_1090, C1 => n_1089, C2 => n_1146, ZN => n_1093);
  g89222 : AOI22D0BWP7T port map(A1 => n_1081, A2 => n_1087, B1 => n_871, B2 => n_1086, ZN => n_1088);
  g89145 : ND4D0BWP7T port map(A1 => n_971, A2 => n_1084, A3 => n_1083, A4 => n_1215, ZN => n_1085);
  g89225 : AOI22D0BWP7T port map(A1 => n_1081, A2 => n_1017, B1 => n_959, B2 => n_1080, ZN => n_1082);
  g89220 : OAI211D1BWP7T port map(A1 => n_1009, A2 => n_857, B => n_981, C => n_703, ZN => n_1079);
  g89177 : ND3D0BWP7T port map(A1 => n_1016, A2 => n_508, A3 => n_836, ZN => n_1078);
  g89178 : IND4D0BWP7T port map(A1 => n_1024, B1 => n_1224, B2 => n_1076, B3 => n_989, ZN => n_1077);
  g89181 : IINR4D0BWP7T port map(A1 => n_1074, A2 => n_1073, B1 => n_986, B2 => n_1072, ZN => n_1075);
  g89218 : ND4D0BWP7T port map(A1 => n_968, A2 => n_768, A3 => n_612, A4 => n_593, ZN => n_1071);
  g89189 : NR4D0BWP7T port map(A1 => n_987, A2 => n_954, A3 => n_953, A4 => n_952, ZN => n_1070);
  g89191 : ND4D0BWP7T port map(A1 => n_993, A2 => n_816, A3 => n_872, A4 => n_1258, ZN => n_1069);
  g89128 : ND4D0BWP7T port map(A1 => n_973, A2 => n_779, A3 => n_1224, A4 => n_1232, ZN => n_1068);
  g89201 : NR4D0BWP7T port map(A1 => n_875, A2 => n_978, A3 => n_1066, A4 => n_647, ZN => n_1067);
  g89186 : IND4D0BWP7T port map(A1 => n_1064, B1 => n_1063, B2 => n_1062, B3 => n_924, ZN => n_1065);
  g89206 : AOI211XD0BWP7T port map(A1 => n_1150, A2 => MISO_shift(66), B => n_990, C => n_705, ZN => n_1061);
  g89208 : OAI221D0BWP7T port map(A1 => n_642, A2 => n_437, B1 => n_896, B2 => n_904, C => n_1019, ZN => n_1060);
  MISO_shift_reg_41 : DFQD1BWP7T port map(CP => clk, D => n_1004, Q => MISO_shift(41));
  g89124 : ND4D0BWP7T port map(A1 => n_947, A2 => n_690, A3 => n_957, A4 => n_1050, ZN => n_1059);
  g89242 : AO222D0BWP7T port map(A1 => n_1026, A2 => n_967, B1 => n_772, B2 => n_1090, C1 => n_681, C2 => n_285, Z => n_1058);
  g89248 : OAI211D1BWP7T port map(A1 => n_1013, A2 => n_392, B => n_944, C => n_133, ZN => n_1057);
  g89165 : IND4D0BWP7T port map(A1 => n_1055, B1 => n_1203, B2 => n_1054, B3 => n_940, ZN => n_1056);
  g89230 : OAI221D0BWP7T port map(A1 => n_1012, A2 => n_1052, B1 => n_704, B2 => n_665, C => n_766, ZN => n_1053);
  g89277 : AOI222D0BWP7T port map(A1 => n_994, A2 => n_1090, B1 => n_870, B2 => n_755, C1 => n_619, C2 => n_1086, ZN => n_1049);
  g89179 : NR4D0BWP7T port map(A1 => n_948, A2 => n_1047, A3 => n_722, A4 => n_1046, ZN => n_1048);
  g89266 : INVD0BWP7T port map(I => n_1045, ZN => n_1147);
  g89187 : IND4D0BWP7T port map(A1 => n_966, B1 => n_1043, B2 => n_1042, B3 => n_776, ZN => n_1044);
  g89192 : ND3D0BWP7T port map(A1 => n_991, A2 => n_1040, A3 => n_1039, ZN => n_1041);
  g89196 : NR4D0BWP7T port map(A1 => n_950, A2 => n_1037, A3 => n_1036, A4 => n_1035, ZN => n_1038);
  g89197 : INR4D0BWP7T port map(A1 => n_1033, B1 => n_1032, B2 => n_1031, B3 => n_920, ZN => n_1034);
  g89198 : NR4D0BWP7T port map(A1 => n_946, A2 => n_1029, A3 => n_1028, A4 => n_409, ZN => n_1030);
  g89199 : AOI211XD0BWP7T port map(A1 => n_1026, A2 => n_992, B => n_960, C => n_786, ZN => n_1027);
  g89188 : IND4D0BWP7T port map(A1 => n_1024, B1 => n_912, B2 => n_788, B3 => n_943, ZN => n_1025);
  MISO_shift_reg_71 : DFQD1BWP7T port map(CP => clk, D => n_976, Q => MISO_shift(71));
  MISO_shift_reg_62 : DFQD1BWP7T port map(CP => clk, D => n_982, Q => MISO_shift(62));
  g89244 : AOI221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(17), B1 => n_721, B2 => n_1092, C => n_906, ZN => n_1023);
  g89234 : ND4D0BWP7T port map(A1 => n_907, A2 => n_682, A3 => n_645, A4 => n_362, ZN => n_1021);
  g89235 : AOI22D0BWP7T port map(A1 => n_1018, A2 => n_1087, B1 => n_841, B2 => n_1146, ZN => n_1020);
  g89241 : AOI22D0BWP7T port map(A1 => n_1018, A2 => n_1017, B1 => n_1150, B2 => MISO_shift(34), ZN => n_1019);
  g89219 : AOI221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(25), B1 => n_795, B2 => n_1015, C => n_925, ZN => n_1016);
  g89273 : OAI32D1BWP7T port map(A1 => n_679, A2 => n_985, A3 => n_139, B1 => n_1013, B2 => n_1012, ZN => n_1014);
  g89275 : OAI222D0BWP7T port map(A1 => n_977, A2 => n_1010, B1 => n_618, B2 => n_853, C1 => n_1009, C2 => n_866, ZN => n_1011);
  g89282 : MAOI22D0BWP7T port map(A1 => n_760, A2 => n_1015, B1 => n_1012, B2 => n_1117, ZN => n_1008);
  g89211 : ND4D0BWP7T port map(A1 => n_917, A2 => n_859, A3 => n_421, A4 => n_277, ZN => n_1007);
  g89190 : NR4D0BWP7T port map(A1 => n_921, A2 => n_887, A3 => n_927, A4 => n_926, ZN => n_1006);
  g89203 : AOI211XD0BWP7T port map(A1 => n_741, A2 => n_941, B => n_929, C => n_739, ZN => n_1005);
  g89209 : IND3D0BWP7T port map(A1 => n_1003, B1 => n_1203, B2 => n_928, ZN => n_1004);
  g89217 : IND4D0BWP7T port map(A1 => n_1001, B1 => n_687, B2 => n_1000, B3 => n_902, ZN => n_1002);
  g89214 : AN3D0BWP7T port map(A1 => n_955, A2 => n_998, A3 => n_997, Z => n_999);
  g89215 : OAI221D0BWP7T port map(A1 => n_995, A2 => n_1010, B1 => n_844, B2 => n_933, C => n_744, ZN => n_996);
  g89287 : AOI211XD0BWP7T port map(A1 => n_706, A2 => full_map_2_2(0), B => n_994, C => n_736, ZN => n_1045);
  g89270 : AOI22D0BWP7T port map(A1 => n_980, A2 => n_992, B1 => n_979, B2 => n_1090, ZN => n_993);
  g89229 : NR3D0BWP7T port map(A1 => n_817, A2 => n_863, A3 => n_425, ZN => n_991);
  g89237 : OAI221D0BWP7T port map(A1 => n_838, A2 => n_1052, B1 => n_1013, B2 => n_370, C => n_913, ZN => n_990);
  g89243 : AN4D0BWP7T port map(A1 => n_988, A2 => n_861, A3 => n_350, A4 => n_347, Z => n_989);
  g89256 : ND4D0BWP7T port map(A1 => n_745, A2 => n_888, A3 => n_471, A4 => n_676, ZN => n_987);
  g89227 : OAI221D0BWP7T port map(A1 => n_945, A2 => n_985, B1 => n_1010, B2 => n_881, C => n_756, ZN => n_986);
  g89264 : IND2D1BWP7T port map(A1 => n_1026, B1 => n_910, ZN => n_1081);
  g89262 : AOI31D0BWP7T port map(A1 => n_635, A2 => n_458, A3 => full_map_9_14(0), B => n_903, ZN => n_1062);
  g89212 : IND4D0BWP7T port map(A1 => n_972, B1 => n_1232, B2 => n_1224, B3 => n_780, ZN => n_982);
  g89276 : AOI22D0BWP7T port map(A1 => n_980, A2 => n_1017, B1 => n_979, B2 => n_1146, ZN => n_981);
  g89279 : OAI22D0BWP7T port map(A1 => n_977, A2 => n_1052, B1 => n_763, B2 => n_833, ZN => n_978);
  g89183 : ND4D0BWP7T port map(A1 => n_892, A2 => n_975, A3 => n_974, A4 => n_1224, ZN => n_976);
  g89185 : NR4D0BWP7T port map(A1 => n_877, A2 => n_972, A3 => n_794, A4 => n_778, ZN => n_973);
  g89200 : NR4D0BWP7T port map(A1 => n_874, A2 => n_970, A3 => n_860, A4 => n_969, ZN => n_971);
  g89272 : AOI32D1BWP7T port map(A1 => n_908, A2 => n_1090, A3 => full_map_5_2(0), B1 => n_980, B2 => n_967, ZN => n_968);
  MISO_shift_reg_18 : DFQD1BWP7T port map(CP => clk, D => n_932, Q => MISO_shift(18));
  MISO_shift_reg_21 : DFQD1BWP7T port map(CP => clk, D => n_919, Q => MISO_shift(21));
  g89254 : OAI221D0BWP7T port map(A1 => n_905, A2 => n_965, B1 => n_1013, B2 => n_521, C => n_502, ZN => n_966);
  g89236 : AOI221D0BWP7T port map(A1 => n_961, A2 => n_1146, B1 => n_1022, B2 => MISO_shift(22), C => n_652, ZN => n_964);
  g89238 : AOI221D0BWP7T port map(A1 => n_962, A2 => n_1080, B1 => n_961, B2 => n_1090, C => n_845, ZN => n_963);
  g89240 : AO211D0BWP7T port map(A1 => n_959, A2 => n_1092, B => n_849, C => n_592, Z => n_960);
  g89228 : INR4D0BWP7T port map(A1 => n_957, B1 => n_847, B2 => n_693, B3 => n_956, ZN => n_958);
  g89246 : NR4D0BWP7T port map(A1 => n_954, A2 => n_832, A3 => n_953, A4 => n_952, ZN => n_955);
  g89251 : AO221D0BWP7T port map(A1 => n_867, A2 => n_1080, B1 => n_1150, B2 => MISO_shift(52), C => n_880, Z => n_951);
  g89252 : ND3D0BWP7T port map(A1 => n_884, A2 => n_842, A3 => n_949, ZN => n_950);
  g89233 : OAI221D0BWP7T port map(A1 => n_862, A2 => n_1013, B1 => n_1010, B2 => n_915, C => n_522, ZN => n_948);
  MISO_shift_reg_36 : DFQD1BWP7T port map(CP => clk, D => n_858, Q => MISO_shift(36));
  g89261 : AOI221D0BWP7T port map(A1 => n_517, A2 => full_map_2_0(0), B1 => n_633, B2 => n_804, C => n_818, ZN => n_1094);
  g89176 : NR4D0BWP7T port map(A1 => n_848, A2 => n_692, A3 => n_691, A4 => n_377, ZN => n_947);
  g89280 : MOAI22D0BWP7T port map(A1 => n_945, A2 => n_901, B1 => n_1022, B2 => MISO_shift(47), ZN => n_946);
  g89295 : OA221D0BWP7T port map(A1 => n_581, A2 => n_1117, B1 => n_373, B2 => n_793, C => n_839, Z => n_944);
  g89271 : AOI222D0BWP7T port map(A1 => n_942, A2 => n_1092, B1 => n_610, B2 => n_941, C1 => n_1150, C2 => MISO_shift(63), ZN => n_943);
  g89210 : NR4D0BWP7T port map(A1 => n_837, A2 => n_939, A3 => n_938, A4 => n_937, ZN => n_940);
  g89353 : INVD0BWP7T port map(I => n_1012, ZN => n_936);
  MISO_shift_reg_63 : DFQD1BWP7T port map(CP => clk, D => n_865, Q => MISO_shift(63));
  g89335 : AOI22D0BWP7T port map(A1 => n_897, A2 => n_1146, B1 => n_935, B2 => MOSI_shift(1), ZN => n_1033);
  MISO_shift_reg_60 : DFQD1BWP7T port map(CP => clk, D => n_864, Q => MISO_shift(60));
  g89349 : AOI22D0BWP7T port map(A1 => n_935, A2 => n_909, B1 => n_574, B2 => n_916, ZN => n_1217);
  g89285 : OAI22D0BWP7T port map(A1 => n_807, A2 => MOSI_shift(1), B1 => n_428, B2 => n_831, ZN => n_983);
  g89267 : MAOI22D0BWP7T port map(A1 => n_961, A2 => n_1080, B1 => n_933, B2 => n_1009, ZN => n_934);
  g89371 : OAI211D1BWP7T port map(A1 => n_893, A2 => n_565, B => n_790, C => n_1258, ZN => n_932);
  g89298 : AOI221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(31), B1 => n_694, B2 => n_941, C => n_784, ZN => n_930);
  g89239 : OAI211D1BWP7T port map(A1 => n_1052, A2 => n_886, B => n_759, C => n_443, ZN => n_929);
  g89247 : NR4D0BWP7T port map(A1 => n_764, A2 => n_775, A3 => n_927, A4 => n_926, ZN => n_928);
  g89253 : OAI221D0BWP7T port map(A1 => n_834, A2 => n_1010, B1 => n_1009, B2 => n_765, C => n_819, ZN => n_925);
  g89255 : AN4D0BWP7T port map(A1 => n_733, A2 => n_923, A3 => n_770, A4 => n_922, Z => n_924);
  g89258 : ND3D0BWP7T port map(A1 => n_796, A2 => n_761, A3 => n_227, ZN => n_921);
  g89259 : OAI211D0BWP7T port map(A1 => n_1117, A2 => n_854, B => n_754, C => n_132, ZN => n_920);
  g89368 : AO211D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(21), B => n_792, C => n_918, Z => n_919);
  g89269 : MAOI22D0BWP7T port map(A1 => n_328, A2 => n_916, B1 => n_915, B2 => n_1117, ZN => n_917);
  g89278 : AOI22D0BWP7T port map(A1 => n_942, A2 => n_1080, B1 => n_876, B2 => n_1146, ZN => n_914);
  g89281 : AOI22D0BWP7T port map(A1 => n_942, A2 => n_1090, B1 => n_718, B2 => n_967, ZN => n_913);
  g89289 : AOI211XD0BWP7T port map(A1 => n_911, A2 => n_1015, B => n_789, C => n_590, ZN => n_912);
  g89302 : ND2D1BWP7T port map(A1 => n_945, A2 => n_910, ZN => n_1018);
  g89284 : AOI22D0BWP7T port map(A1 => n_806, A2 => MOSI_shift(1), B1 => n_800, B2 => n_909, ZN => n_1040);
  MISO_shift_reg_42 : DFQD1BWP7T port map(CP => clk, D => n_823, Q => MISO_shift(42));
  g89382 : AOI211XD0BWP7T port map(A1 => n_908, A2 => full_map_2_2(0), B => n_777, C => n_767, ZN => n_1012);
  g89328 : AOI22D0BWP7T port map(A1 => n_899, A2 => n_1080, B1 => n_898, B2 => n_1087, ZN => n_907);
  g89324 : OAI22D0BWP7T port map(A1 => n_905, A2 => n_985, B1 => n_904, B2 => n_827, ZN => n_906);
  g89323 : OAI32D0BWP7T port map(A1 => n_519, A2 => n_455, A3 => n_42, B1 => MOSI_shift(1), B2 => n_894, ZN => n_903);
  g89330 : MAOI22D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(13), B1 => n_905, B2 => n_901, ZN => n_902);
  g89331 : AOI22D0BWP7T port map(A1 => n_899, A2 => n_1146, B1 => n_898, B2 => n_1017, ZN => n_900);
  MISO_shift_reg_54 : DFQD1BWP7T port map(CP => clk, D => n_813, Q => MISO_shift(54));
  MISO_shift_reg_27 : DFQD1BWP7T port map(CP => clk, D => n_852, Q => MISO_shift(27));
  MISO_shift_reg_57 : DFQD1BWP7T port map(CP => clk, D => n_808, Q => MISO_shift(57));
  MISO_shift_reg_24 : DFQD1BWP7T port map(CP => clk, D => n_810, Q => MISO_shift(24));
  g89354 : INVD0BWP7T port map(I => n_977, ZN => n_994);
  MISO_shift_reg_69 : DFQD1BWP7T port map(CP => clk, D => n_815, Q => MISO_shift(69));
  MISO_shift_reg_39 : DFQD1BWP7T port map(CP => clk, D => n_809, Q => MISO_shift(39));
  MISO_shift_reg_66 : DFQD1BWP7T port map(CP => clk, D => n_811, Q => MISO_shift(66));
  MISO_shift_reg_51 : DFQD1BWP7T port map(CP => clk, D => n_805, Q => MISO_shift(51));
  g89339 : MAOI22D0BWP7T port map(A1 => n_897, A2 => n_1080, B1 => n_896, B2 => n_829, ZN => n_1076);
  g89341 : OAI22D0BWP7T port map(A1 => n_895, A2 => n_901, B1 => n_729, B2 => n_896, ZN => n_1047);
  g89346 : OAI22D0BWP7T port map(A1 => n_895, A2 => n_909, B1 => n_713, B2 => n_604, ZN => n_1113);
  g89348 : OAI22D0BWP7T port map(A1 => n_856, A2 => n_901, B1 => n_894, B2 => n_893, ZN => n_1003);
  g89319 : IOA21D1BWP7T port map(A1 => n_641, A2 => full_map_2_2(0), B => n_945, ZN => n_1026);
  g89249 : NR4D0BWP7T port map(A1 => n_891, A2 => n_609, A3 => n_890, A4 => n_889, ZN => n_892);
  g89374 : AOI221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(58), B1 => n_1150, B2 => MISO_shift(57), C => n_725, ZN => n_888);
  g89300 : OAI221D0BWP7T port map(A1 => n_886, A2 => n_1013, B1 => n_985, B2 => n_843, C => n_742, ZN => n_887);
  g89299 : AOI221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(37), B1 => n_1150, B2 => MISO_shift(36), C => n_746, ZN => n_885);
  g89397 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(29), B1 => n_883, B2 => n_893, ZN => n_884);
  g89405 : MOAI22D0BWP7T port map(A1 => n_881, A2 => n_1013, B1 => n_1022, B2 => MISO_shift(35), ZN => n_882);
  g89408 : MOAI22D0BWP7T port map(A1 => n_881, A2 => n_1117, B1 => n_1022, B2 => MISO_shift(53), ZN => n_880);
  g89373 : AOI221D0BWP7T port map(A1 => n_878, A2 => n_967, B1 => n_723, B2 => n_1086, C => n_714, ZN => n_879);
  g89250 : AO221D0BWP7T port map(A1 => n_787, A2 => n_967, B1 => n_876, B2 => n_1092, C => n_753, Z => n_877);
  g89257 : OAI211D1BWP7T port map(A1 => n_1117, A2 => n_873, B => n_720, C => n_237, ZN => n_875);
  g89268 : OAI221D0BWP7T port map(A1 => n_873, A2 => n_1013, B1 => n_589, B2 => n_904, C => n_677, ZN => n_874);
  g89291 : AOI221D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(15), B1 => n_871, B2 => n_941, C => n_735, ZN => n_872);
  g89286 : OAI222D0BWP7T port map(A1 => n_873, A2 => n_965, B1 => MOSI_shift(5), B2 => n_494, C1 => n_801, C2 => n_638, ZN => n_1155);
  g89381 : IOA21D1BWP7T port map(A1 => n_855, A2 => full_map_2_2(0), B => n_905, ZN => n_980);
  g89385 : AOI221D0BWP7T port map(A1 => n_870, A2 => full_map_2_14(0), B1 => n_869, B2 => n_555, C => n_824, ZN => n_977);
  g89334 : MAOI22D0BWP7T port map(A1 => n_867, A2 => n_1146, B1 => n_866, B2 => n_1010, ZN => n_868);
  g89360 : OAI221D0BWP7T port map(A1 => n_812, A2 => n_901, B1 => n_985, B2 => n_683, C => n_717, ZN => n_865);
  g89355 : OAI221D0BWP7T port map(A1 => n_814, A2 => n_1052, B1 => n_851, B2 => n_545, C => n_234, ZN => n_864);
  g89320 : OAI22D0BWP7T port map(A1 => n_862, A2 => n_1117, B1 => n_448, B2 => n_1010, ZN => n_863);
  g89325 : AOI32D1BWP7T port map(A1 => n_825, A2 => n_992, A3 => full_map_1_13(1), B1 => n_867, B2 => n_1092, ZN => n_861);
  g89327 : OAI21D0BWP7T port map(A1 => n_862, A2 => n_1010, B => n_438, ZN => n_860);
  g89332 : MAOI22D0BWP7T port map(A1 => n_556, A2 => n_345, B1 => n_862, B2 => n_1052, ZN => n_859);
  g89301 : IND3D1BWP7T port map(A1 => n_585, B1 => n_399, B2 => n_731, ZN => n_858);
  g89303 : AN2D0BWP7T port map(A1 => n_915, A2 => n_857, Z => n_995);
  g89340 : OAI22D0BWP7T port map(A1 => n_856, A2 => n_909, B1 => n_528, B2 => MOSI_shift(8), ZN => n_1064);
  g89344 : AOI222D0BWP7T port map(A1 => n_828, A2 => n_967, B1 => n_119, B2 => n_749, C1 => n_750, C2 => n_1087, ZN => n_988);
  g89345 : AOI22D0BWP7T port map(A1 => n_867, A2 => n_1017, B1 => n_855, B2 => n_670, ZN => n_1129);
  g89337 : OAI222D0BWP7T port map(A1 => n_854, A2 => n_985, B1 => n_965, B2 => n_830, C1 => n_751, C2 => n_826, ZN => n_972);
  g89315 : OA21D0BWP7T port map(A1 => n_856, A2 => n_893, B => n_1215, Z => n_1054);
  g89338 : OAI222D0BWP7T port map(A1 => n_873, A2 => n_985, B1 => n_664, B2 => n_667, C1 => n_32, C2 => n_853, ZN => n_1193);
  g89369 : OAI221D0BWP7T port map(A1 => n_822, A2 => n_1052, B1 => n_851, B2 => n_605, C => n_267, ZN => n_852);
  g89370 : AOI211D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(4), B => n_680, C => n_509, ZN => n_850);
  g89292 : OAI221D0BWP7T port map(A1 => n_375, A2 => n_651, B1 => n_710, B2 => n_853, C => n_737, ZN => n_849);
  g89232 : IND4D0BWP7T port map(A1 => n_847, B1 => n_846, B2 => n_696, B3 => n_659, ZN => n_848);
  g89401 : OAI22D0BWP7T port map(A1 => n_886, A2 => n_844, B1 => n_843, B2 => n_901, ZN => n_845);
  g89403 : AOI22D0BWP7T port map(A1 => n_841, A2 => n_1080, B1 => n_1150, B2 => MISO_shift(28), ZN => n_842);
  g89407 : AOI22D0BWP7T port map(A1 => n_959, A2 => n_1090, B1 => n_1150, B2 => MISO_shift(51), ZN => n_840);
  g89409 : MAOI22D0BWP7T port map(A1 => n_341, A2 => n_820, B1 => n_838, B2 => n_1010, ZN => n_839);
  g89290 : IND4D0BWP7T port map(A1 => n_653, B1 => n_430, B2 => n_346, B3 => n_836, ZN => n_837);
  g89245 : OAI221D0BWP7T port map(A1 => n_834, A2 => n_833, B1 => n_1117, B2 => n_678, C => n_643, ZN => n_835);
  g89422 : CKND2D1BWP7T port map(A1 => n_716, A2 => n_620, ZN => n_832);
  g89283 : OAI222D0BWP7T port map(A1 => n_799, A2 => n_909, B1 => n_831, B2 => n_669, C1 => n_548, C2 => n_802, ZN => n_1178);
  g89415 : OA22D0BWP7T port map(A1 => n_830, A2 => n_1010, B1 => n_578, B2 => n_220, Z => n_975);
  g89440 : OAI21D0BWP7T port map(A1 => n_829, A2 => n_774, B => n_726, ZN => n_935);
  g89260 : AOI211D0BWP7T port map(A1 => n_797, A2 => n_992, B => n_436, C => n_243, ZN => n_1127);
  g89416 : AOI22D0BWP7T port map(A1 => n_752, A2 => n_967, B1 => n_447, B2 => n_1087, ZN => n_1102);
  g89413 : OAI22D0BWP7T port map(A1 => n_747, A2 => n_893, B1 => n_730, B2 => n_771, ZN => n_956);
  g89412 : MAOI22D0BWP7T port map(A1 => n_828, A2 => n_1087, B1 => n_827, B2 => n_829, ZN => n_1181);
  g89417 : OA22D0BWP7T port map(A1 => n_803, A2 => n_1052, B1 => n_826, B2 => n_1224, Z => n_1192);
  g89383 : AOI21D0BWP7T port map(A1 => n_825, A2 => full_map_2_14(0), B => n_824, ZN => n_945);
  g89365 : OAI221D0BWP7T port map(A1 => n_822, A2 => n_1117, B1 => n_1010, B2 => n_791, C => n_624, ZN => n_823);
  g89296 : AOI221D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(21), B1 => n_688, B2 => n_820, C => n_686, ZN => n_821);
  g89297 : AOI221D0BWP7T port map(A1 => n_384, A2 => n_1086, B1 => n_908, B2 => n_526, C => n_701, ZN => n_819);
  g89322 : OAI32D1BWP7T port map(A1 => n_244, A2 => n_965, A3 => n_748, B1 => n_893, B2 => n_773, ZN => n_818);
  g89326 : OAI22D0BWP7T port map(A1 => n_873, A2 => n_1052, B1 => n_762, B2 => n_893, ZN => n_817);
  g89294 : AOI221D0BWP7T port map(A1 => n_855, A2 => n_14, B1 => n_1022, B2 => MISO_shift(16), C => n_702, ZN => n_816);
  g89364 : OAI211D1BWP7T port map(A1 => n_1010, A2 => n_814, B => n_654, C => n_534, ZN => n_815);
  g89363 : OAI211D1BWP7T port map(A1 => n_965, A2 => n_812, B => n_656, C => n_533, ZN => n_813);
  g89361 : OAI211D1BWP7T port map(A1 => n_985, A2 => n_812, B => n_658, C => n_529, ZN => n_811);
  g89359 : OAI211D1BWP7T port map(A1 => n_1013, A2 => n_822, B => n_530, C => n_657, ZN => n_810);
  g89358 : OAI211D1BWP7T port map(A1 => n_1010, A2 => n_822, B => n_536, C => n_650, ZN => n_809);
  g89357 : OAI211D1BWP7T port map(A1 => n_1013, A2 => n_814, B => n_531, C => n_648, ZN => n_808);
  g89352 : INVD0BWP7T port map(I => n_806, ZN => n_807);
  g89356 : OAI211D1BWP7T port map(A1 => n_893, A2 => n_812, B => n_407, C => n_661, ZN => n_805);
  g89336 : AOI21D0BWP7T port map(A1 => n_482, A2 => n_804, B => n_743, ZN => n_1084);
  g89350 : OAI22D0BWP7T port map(A1 => n_873, A2 => n_901, B1 => n_803, B2 => n_1013, ZN => n_1171);
  MISO_shift_reg_45 : DFQD1BWP7T port map(CP => clk, D => n_734, Q => MISO_shift(45));
  g89347 : OAI22D0BWP7T port map(A1 => n_854, A2 => n_893, B1 => n_802, B2 => n_801, ZN => n_1122);
  g89343 : OAI32D1BWP7T port map(A1 => n_798, A2 => n_466, A3 => n_1231, B1 => n_893, B2 => n_873, ZN => n_1111);
  g89342 : MAOI22D0BWP7T port map(A1 => n_800, A2 => MOSI_shift(1), B1 => n_799, B2 => MOSI_shift(1), ZN => n_1160);
  g89351 : MOAI22D0BWP7T port map(A1 => n_583, A2 => n_798, B1 => n_797, B2 => n_1080, ZN => n_1132);
  g89404 : AOI22D0BWP7T port map(A1 => n_613, A2 => n_941, B1 => n_795, B2 => n_1086, ZN => n_796);
  g89372 : OAI221D0BWP7T port map(A1 => n_631, A2 => n_844, B1 => n_793, B2 => n_827, C => n_431, ZN => n_794);
  g89431 : OAI221D0BWP7T port map(A1 => n_563, A2 => n_570, B1 => n_833, B2 => n_791, C => n_644, ZN => n_792);
  g89429 : AOI221D0BWP7T port map(A1 => n_663, A2 => full_map_2_1(2), B1 => n_1150, B2 => MISO_shift(17), C => n_576, ZN => n_790);
  g89427 : NR2D0BWP7T port map(A1 => n_838, A2 => n_1013, ZN => n_789);
  g89426 : AOI221D0BWP7T port map(A1 => n_787, A2 => n_992, B1 => n_1022, B2 => MISO_shift(64), C => n_582, ZN => n_788);
  g89388 : MOAI22D0BWP7T port map(A1 => n_785, A2 => n_1117, B1 => n_787, B2 => n_1087, ZN => n_786);
  g89391 : OAI22D0BWP7T port map(A1 => n_782, A2 => n_833, B1 => n_785, B2 => n_1013, ZN => n_784);
  g89392 : OAI22D0BWP7T port map(A1 => n_782, A2 => n_781, B1 => n_785, B2 => n_1010, ZN => n_783);
  g89367 : IINR4D0BWP7T port map(A1 => n_779, A2 => n_364, B1 => n_623, B2 => n_778, ZN => n_780);
  g89418 : INVD0BWP7T port map(I => n_862, ZN => n_777);
  g89424 : AOI211XD0BWP7T port map(A1 => n_1150, A2 => MISO_shift(4), B => n_577, C => n_459, ZN => n_776);
  g89425 : AO221D0BWP7T port map(A1 => n_769, A2 => n_1080, B1 => n_1150, B2 => MISO_shift(40), C => n_594, Z => n_775);
  g89378 : OAI21D0BWP7T port map(A1 => n_575, A2 => n_774, B => n_773, ZN => n_806);
  g89437 : OR2D1BWP7T port map(A1 => n_841, A2 => n_772, Z => n_899);
  g89379 : IND2D1BWP7T port map(A1 => n_871, B1 => n_873, ZN => n_961);
  g89380 : AOI21D0BWP7T port map(A1 => n_524, A2 => n_118, B => n_797, ZN => n_915);
  g89384 : OAI21D0BWP7T port map(A1 => n_771, A2 => n_468, B => n_854, ZN => n_942);
  g89505 : AOI222D0BWP7T port map(A1 => n_769, A2 => n_1146, B1 => n_758, B2 => full_map_1_13(1), C1 => n_1150, C2 => MISO_shift(43), ZN => n_770);
  g89333 : AOI22D0BWP7T port map(A1 => n_979, A2 => n_1092, B1 => n_767, B2 => n_1086, ZN => n_768);
  g89329 : OA22D0BWP7T port map(A1 => n_834, A2 => n_844, B1 => n_833, B2 => n_765, Z => n_766);
  g89458 : OAI222D0BWP7T port map(A1 => n_763, A2 => n_844, B1 => n_985, B2 => n_762, C1 => n_965, C2 => n_646, ZN => n_764);
  g89459 : AOI22D0BWP7T port map(A1 => n_878, A2 => n_1017, B1 => n_760, B2 => n_820, ZN => n_761);
  g89321 : AOI222D0BWP7T port map(A1 => n_758, A2 => full_map_1_13(0), B1 => n_539, B2 => n_1015, C1 => n_1150, C2 => MISO_shift(42), ZN => n_759);
  g89293 : AOI221D0BWP7T port map(A1 => n_962, A2 => n_820, B1 => n_1022, B2 => MISO_shift(52), C => n_527, ZN => n_757);
  g89493 : AOI221D0BWP7T port map(A1 => n_825, A2 => n_755, B1 => n_1022, B2 => MISO_shift(50), C => n_588, ZN => n_756);
  g89496 : AOI221D0BWP7T port map(A1 => n_363, A2 => n_1080, B1 => n_1150, B2 => MISO_shift(67), C => n_622, ZN => n_754);
  g89288 : OAI211D0BWP7T port map(A1 => n_401, A2 => n_499, B => n_611, C => n_580, ZN => n_753);
  g89445 : AOI21D0BWP7T port map(A1 => n_870, A2 => full_map_0_14(0), B => n_752, ZN => n_894);
  g89487 : OAI21D0BWP7T port map(A1 => n_294, A2 => n_751, B => n_830, ZN => n_897);
  g89476 : AO222D0BWP7T port map(A1 => n_750, A2 => n_909, B1 => n_128, B2 => n_749, C1 => n_217, C2 => n_493, Z => n_1031);
  MISO_shift_reg_15 : DFQD1BWP7T port map(CP => clk, D => n_700, Q => MISO_shift(15));
  MISO_shift_reg_33 : DFQD1BWP7T port map(CP => clk, D => n_699, Q => MISO_shift(33));
  MISO_shift_reg_48 : DFQD1BWP7T port map(CP => clk, D => n_684, Q => MISO_shift(48));
  g89439 : OA21D0BWP7T port map(A1 => n_748, A2 => n_287, B => n_747, Z => n_895);
  g89450 : AOI211XD0BWP7T port map(A1 => n_457, A2 => full_map_2_14(0), B => n_728, C => n_727, ZN => n_905);
  g89411 : MOAI22D0BWP7T port map(A1 => n_738, A2 => n_833, B1 => n_760, B2 => n_1086, ZN => n_746);
  g89387 : AOI32D1BWP7T port map(A1 => n_501, A2 => n_629, A3 => full_map_10_11(0), B1 => n_962, B2 => n_1090, ZN => n_745);
  g89389 : AOI22D0BWP7T port map(A1 => n_1091, A2 => n_1146, B1 => n_1150, B2 => MISO_shift(6), ZN => n_744);
  g89390 : OAI22D0BWP7T port map(A1 => n_673, A2 => n_901, B1 => n_748, B2 => n_390, ZN => n_743);
  g89393 : AOI22D0BWP7T port map(A1 => n_962, A2 => n_1146, B1 => n_741, B2 => n_1015, ZN => n_742);
  g89395 : AOI22D0BWP7T port map(A1 => n_962, A2 => n_1092, B1 => n_1022, B2 => MISO_shift(55), ZN => n_740);
  g89398 : MOAI22D0BWP7T port map(A1 => n_738, A2 => n_1013, B1 => n_760, B2 => n_1092, ZN => n_739);
  g89402 : AOI22D0BWP7T port map(A1 => n_962, A2 => n_1086, B1 => n_736, B2 => n_820, ZN => n_737);
  g89406 : AO22D0BWP7T port map(A1 => n_1091, A2 => n_1092, B1 => n_1080, B2 => n_1089, Z => n_735);
  g89375 : AO221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(45), B1 => n_1150, B2 => MISO_shift(44), C => n_606, Z => n_734);
  g89463 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(44), B1 => n_763, B2 => n_1013, ZN => n_733);
  g89461 : MOAI22D0BWP7T port map(A1 => n_782, A2 => n_844, B1 => n_871, B2 => n_820, ZN => n_732);
  g89457 : AOI222D0BWP7T port map(A1 => n_564, A2 => n_967, B1 => n_1150, B2 => MISO_shift(35), C1 => n_1022, C2 => MISO_shift(36), ZN => n_731);
  g89441 : OAI221D0BWP7T port map(A1 => n_441, A2 => n_662, B1 => n_252, B2 => n_326, C => n_614, ZN => n_824);
  g89414 : OAI222D0BWP7T port map(A1 => n_730, A2 => n_1231, B1 => n_279, B2 => n_729, C1 => n_893, C2 => n_674, ZN => n_970);
  g89447 : AOI211D0BWP7T port map(A1 => n_542, A2 => full_map_0_13(0), B => n_504, C => n_569, ZN => n_856);
  g89419 : INVD1BWP7T port map(I => n_854, ZN => n_867);
  g89451 : NR3D0BWP7T port map(A1 => n_728, A2 => n_727, A3 => n_434, ZN => n_862);
  g89488 : INVD0BWP7T port map(I => n_828, ZN => n_726);
  g89467 : MOAI22D0BWP7T port map(A1 => n_724, A2 => n_1010, B1 => n_723, B2 => n_820, ZN => n_725);
  g89362 : AO221D0BWP7T port map(A1 => n_721, A2 => n_1146, B1 => n_1150, B2 => MISO_shift(7), C => n_584, Z => n_722);
  g89540 : AOI22D0BWP7T port map(A1 => n_769, A2 => n_941, B1 => n_715, B2 => n_1080, ZN => n_720);
  g89539 : AOI22D0BWP7T port map(A1 => n_540, A2 => n_1015, B1 => n_718, B2 => n_1087, ZN => n_719);
  g89498 : AOI222D0BWP7T port map(A1 => n_498, A2 => n_1090, B1 => n_1022, B2 => MISO_shift(63), C1 => n_1150, C2 => MISO_shift(62), ZN => n_717);
  g89495 : AOI222D0BWP7T port map(A1 => n_715, A2 => n_1090, B1 => n_1150, B2 => MISO_shift(58), C1 => n_1022, C2 => MISO_shift(59), ZN => n_716);
  g89466 : MOAI22D0BWP7T port map(A1 => n_724, A2 => n_1009, B1 => n_1150, B2 => MISO_shift(54), ZN => n_714);
  g89486 : AOI22D0BWP7T port map(A1 => n_707, A2 => n_1092, B1 => n_626, B2 => n_1090, ZN => n_1123);
  g89481 : OAI22D0BWP7T port map(A1 => n_712, A2 => n_798, B1 => n_853, B2 => n_672, ZN => n_969);
  g89480 : OAI22D0BWP7T port map(A1 => n_709, A2 => n_711, B1 => n_713, B2 => n_708, ZN => n_1110);
  g89514 : INR2D0BWP7T port map(A1 => n_408, B1 => n_898, ZN => n_883);
  g89470 : OAI22D0BWP7T port map(A1 => n_712, A2 => n_711, B1 => n_748, B2 => n_710, ZN => n_1154);
  g89479 : OAI22D0BWP7T port map(A1 => n_709, A2 => n_798, B1 => n_552, B2 => n_708, ZN => n_1153);
  g89474 : MOAI22D0BWP7T port map(A1 => n_627, A2 => n_666, B1 => n_750, B2 => n_967, ZN => n_891);
  MISO_shift_reg_30 : DFQD1BWP7T port map(CP => clk, D => n_591, Q => MISO_shift(30));
  g89471 : MAOI22D0BWP7T port map(A1 => n_707, A2 => n_1090, B1 => n_802, B2 => n_634, ZN => n_1074);
  g89524 : AOI21D0BWP7T port map(A1 => n_706, A2 => full_map_3_2(1), B => n_587, ZN => n_881);
  g89433 : OAI221D0BWP7T port map(A1 => n_599, A2 => n_616, B1 => n_704, B2 => n_632, C => n_541, ZN => n_705);
  g89399 : MAOI22D0BWP7T port map(A1 => n_767, A2 => n_941, B1 => n_933, B2 => n_833, ZN => n_703);
  g89400 : MOAI22D0BWP7T port map(A1 => n_933, A2 => n_781, B1 => n_767, B2 => n_820, ZN => n_702);
  g89410 : OAI22D0BWP7T port map(A1 => n_933, A2 => n_1117, B1 => n_843, B2 => n_965, ZN => n_701);
  g89421 : OAI221D0BWP7T port map(A1 => n_698, A2 => n_893, B1 => n_1013, B2 => n_697, C => n_228, ZN => n_700);
  g89423 : OAI221D0BWP7T port map(A1 => n_698, A2 => n_901, B1 => n_1010, B2 => n_697, C => n_232, ZN => n_699);
  g89428 : AOI221D0BWP7T port map(A1 => n_660, A2 => full_map_3_5(0), B1 => n_640, B2 => n_675, C => n_342, ZN => n_696);
  g89430 : AO221D0BWP7T port map(A1 => n_694, A2 => n_820, B1 => n_1022, B2 => MISO_shift(46), C => n_424, Z => n_695);
  g89432 : IIND4D0BWP7T port map(A1 => n_692, A2 => n_691, B1 => n_690, B2 => n_311, ZN => n_693);
  g89396 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1086, B1 => n_1022, B2 => MISO_shift(19), ZN => n_689);
  g89434 : AOI31D0BWP7T port map(A1 => n_855, A2 => n_992, A3 => full_map_3_2(1), B => n_535, ZN => n_687);
  g89394 : OAI22D0BWP7T port map(A1 => n_933, A2 => n_1010, B1 => n_765, B2 => n_781, ZN => n_686);
  g89386 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(10), B1 => n_933, B2 => n_1013, ZN => n_685);
  g89497 : OAI211D1BWP7T port map(A1 => n_893, A2 => n_683, B => n_476, C => n_176, ZN => n_684);
  g89455 : AOI22D0BWP7T port map(A1 => n_571, A2 => n_941, B1 => n_681, B2 => n_601, ZN => n_682);
  g89460 : OAI32D1BWP7T port map(A1 => n_679, A2 => n_343, A3 => n_348, B1 => n_1010, B2 => n_678, ZN => n_680);
  g89462 : AOI22D0BWP7T port map(A1 => n_721, A2 => n_1090, B1 => n_1022, B2 => MISO_shift(20), ZN => n_677);
  g89464 : AOI22D0BWP7T port map(A1 => n_741, A2 => n_1086, B1 => n_870, B2 => n_675, ZN => n_676);
  g89435 : OAI211D1BWP7T port map(A1 => n_628, A2 => n_729, B => n_674, C => n_483, ZN => n_800);
  g89442 : OA21D0BWP7T port map(A1 => n_748, A2 => n_304, B => n_673, Z => n_773);
  g89484 : OAI22D0BWP7T port map(A1 => n_671, A2 => n_711, B1 => n_625, B2 => n_798, ZN => n_1121);
  g89468 : OAI22D0BWP7T port map(A1 => n_472, A2 => n_901, B1 => n_639, B2 => n_672, ZN => n_939);
  g89469 : OAI22D0BWP7T port map(A1 => n_671, A2 => n_798, B1 => n_910, B2 => n_637, ZN => n_1072);
  g89472 : MOAI22D0BWP7T port map(A1 => n_668, A2 => n_798, B1 => n_908, B2 => n_670, ZN => n_1177);
  g89473 : OAI22D0BWP7T port map(A1 => n_470, A2 => n_1010, B1 => n_771, B2 => n_909, ZN => n_1131);
  g89475 : OAI22D0BWP7T port map(A1 => n_910, A2 => MOSI_shift(5), B1 => n_669, B2 => n_708, ZN => n_1029);
  g89477 : OAI22D0BWP7T port map(A1 => n_668, A2 => n_711, B1 => n_667, B2 => n_666, ZN => n_1182);
  g89482 : OAI22D0BWP7T port map(A1 => n_668, A2 => n_1052, B1 => n_665, B2 => n_664, ZN => n_1066);
  g89483 : AOI22D0BWP7T port map(A1 => n_442, A2 => MOSI_shift(2), B1 => n_663, B2 => full_map_4_0(0), ZN => n_949);
  g89446 : OAI211D1BWP7T port map(A1 => n_662, A2 => n_109, B => n_410, C => n_479, ZN => n_797);
  g89452 : AOI221D0BWP7T port map(A1 => n_630, A2 => full_map_14_13(0), B1 => n_505, B2 => full_map_14_11(0), C => n_475, ZN => n_854);
  g89453 : AOI211XD0BWP7T port map(A1 => n_484, A2 => full_map_14_1(0), B => n_445, C => n_495, ZN => n_873);
  g89549 : AOI22D0BWP7T port map(A1 => n_660, A2 => full_map_4_1(2), B1 => n_1150, B2 => MISO_shift(50), ZN => n_661);
  g89366 : AOI211D0BWP7T port map(A1 => n_344, A2 => n_385, B => n_477, C => n_327, ZN => n_659);
  g89566 : AOI22D0BWP7T port map(A1 => n_655, A2 => n_1092, B1 => n_1150, B2 => MISO_shift(65), ZN => n_658);
  g89563 : AOI22D0BWP7T port map(A1 => n_649, A2 => n_1146, B1 => n_1150, B2 => MISO_shift(23), ZN => n_657);
  g89560 : AOI22D0BWP7T port map(A1 => n_655, A2 => n_1080, B1 => n_1150, B2 => MISO_shift(53), ZN => n_656);
  g89559 : AOI22D0BWP7T port map(A1 => n_655, A2 => n_1090, B1 => n_1150, B2 => MISO_shift(68), ZN => n_654);
  g89557 : MOAI22D0BWP7T port map(A1 => n_762, A2 => n_965, B1 => n_597, B2 => n_1092, ZN => n_653);
  g89556 : OAI22D0BWP7T port map(A1 => n_665, A2 => n_651, B1 => n_843, B2 => n_893, ZN => n_652);
  g89554 : AOI22D0BWP7T port map(A1 => n_649, A2 => n_1090, B1 => n_1150, B2 => MISO_shift(38), ZN => n_650);
  g89553 : AOI22D0BWP7T port map(A1 => n_660, A2 => full_map_2_1(2), B1 => n_1022, B2 => MISO_shift(57), ZN => n_648);
  g89552 : OAI22D0BWP7T port map(A1 => n_762, A2 => n_901, B1 => n_646, B2 => n_893, ZN => n_647);
  g89548 : AOI22D0BWP7T port map(A1 => n_660, A2 => full_map_6_2(0), B1 => n_1150, B2 => MISO_shift(27), ZN => n_645);
  g89545 : AOI22D0BWP7T port map(A1 => n_649, A2 => n_1080, B1 => n_1150, B2 => MISO_shift(20), ZN => n_644);
  g89543 : AOI22D0BWP7T port map(A1 => n_663, A2 => full_map_1_2(0), B1 => n_1022, B2 => MISO_shift(7), ZN => n_643);
  g89515 : OA221D0BWP7T port map(A1 => n_642, A2 => n_598, B1 => n_36, B2 => n_537, C => n_332, Z => n_1143);
  g89507 : INR2D1BWP7T port map(A1 => n_671, B1 => n_707, ZN => n_803);
  g89508 : OAI222D0BWP7T port map(A1 => n_669, A2 => n_603, B1 => n_1010, B2 => n_547, C1 => n_419, C2 => n_802, ZN => n_954);
  g89509 : AOI221D0BWP7T port map(A1 => n_641, A2 => full_map_0_5(0), B1 => n_640, B2 => full_map_0_13(0), C => n_463, ZN => n_747);
  g89601 : OAI32D1BWP7T port map(A1 => full_map_6_0(0), A2 => n_798, A3 => n_639, B1 => n_558, B2 => n_638, ZN => n_1001);
  g89580 : MAOI22D0BWP7T port map(A1 => n_518, A2 => n_512, B1 => n_636, B2 => n_637, ZN => n_1208);
  g89520 : OAI32D1BWP7T port map(A1 => n_554, A2 => n_1117, A3 => n_771, B1 => MOSI_shift(5), B2 => n_636, ZN => n_1109);
  g89518 : AOI31D0BWP7T port map(A1 => n_635, A2 => n_596, A3 => full_map_5_14(0), B => n_562, ZN => n_923);
  g89579 : OAI32D1BWP7T port map(A1 => n_366, A2 => n_634, A3 => n_1224, B1 => n_985, B2 => n_573, ZN => n_1028);
  g89513 : AO221D0BWP7T port map(A1 => n_633, A2 => n_489, B1 => n_706, B2 => full_map_0_2(0), C => n_544, Z => n_752);
  g89528 : OA21D0BWP7T port map(A1 => n_632, A2 => n_579, B => n_631, Z => n_838);
  g89525 : IND2D1BWP7T port map(A1 => n_694, B1 => n_586, ZN => n_959);
  g89618 : AOI21D0BWP7T port map(A1 => n_706, A2 => full_map_1_1(2), B => n_718, ZN => n_814);
  g89530 : INR2XD0BWP7T port map(A1 => n_724, B1 => n_769, ZN => n_886);
  g89526 : AOI221D0BWP7T port map(A1 => n_630, A2 => full_map_14_12(0), B1 => n_124, B2 => n_629, C => n_507, ZN => n_830);
  g89527 : OAI221D0BWP7T port map(A1 => n_568, A2 => n_628, B1 => n_566, B2 => n_627, C => n_525, ZN => n_828);
  g89523 : IND2D1BWP7T port map(A1 => n_626, B1 => n_625, ZN => n_841);
  g89628 : AOI21D0BWP7T port map(A1 => n_641, A2 => full_map_1_1(2), B => n_787, ZN => n_812);
  g89499 : AOI222D0BWP7T port map(A1 => n_380, A2 => n_1086, B1 => n_1022, B2 => MISO_shift(42), C1 => n_1150, C2 => MISO_shift(41), ZN => n_624);
  g89690 : MOAI22D0BWP7T port map(A1 => n_853, A2 => n_621, B1 => n_360, B2 => n_1080, ZN => n_623);
  g89691 : MOAI22D0BWP7T port map(A1 => n_639, A2 => n_621, B1 => n_1022, B2 => MISO_shift(68), ZN => n_622);
  g89695 : MAOI22D0BWP7T port map(A1 => n_619, A2 => n_820, B1 => n_639, B2 => n_618, ZN => n_620);
  g89688 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(70), B1 => n_669, B2 => n_616, ZN => n_617);
  g89492 : AOI32D0BWP7T port map(A1 => n_641, A2 => n_1017, A3 => full_map_4_2(0), B1 => n_694, B2 => n_1015, ZN => n_615);
  g89490 : AOI222D0BWP7T port map(A1 => n_630, A2 => full_map_14_14(0), B1 => n_351, B2 => n_629, C1 => n_480, C2 => full_map_14_2(0), ZN => n_614);
  g89489 : INVD0BWP7T port map(I => n_738, ZN => n_613);
  g89465 : AOI22D0BWP7T port map(A1 => n_549, A2 => n_820, B1 => n_1022, B2 => MISO_shift(13), ZN => n_612);
  g89456 : AOI222D0BWP7T port map(A1 => n_610, A2 => n_1015, B1 => n_1022, B2 => MISO_shift(61), C1 => n_174, C2 => n_1146, ZN => n_611);
  g89420 : IND3D0BWP7T port map(A1 => n_608, B1 => n_361, B2 => n_607, ZN => n_609);
  g89454 : OAI221D0BWP7T port map(A1 => n_605, A2 => n_45, B1 => n_1117, B2 => n_791, C => n_423, ZN => n_606);
  g89485 : OAI32D1BWP7T port map(A1 => full_map_6_0(0), A2 => n_1052, A3 => n_665, B1 => n_439, B2 => n_444, ZN => n_1036);
  g89698 : OAI22D0BWP7T port map(A1 => n_400, A2 => n_604, B1 => n_713, B2 => n_831, ZN => n_1139);
  g89436 : AOI221D0BWP7T port map(A1 => n_825, A2 => full_map_0_14(0), B1 => n_600, B2 => n_523, C => n_602, ZN => n_799);
  g89719 : MOAI22D0BWP7T port map(A1 => n_642, A2 => n_603, B1 => n_520, B2 => n_1146, ZN => n_927);
  g89478 : AO22D0BWP7T port map(A1 => n_602, A2 => n_967, B1 => n_601, B2 => n_600, Z => n_1100);
  g89701 : OAI22D0BWP7T port map(A1 => n_599, A2 => n_550, B1 => n_84, B2 => n_513, ZN => n_1035);
  g89709 : OAI22D0BWP7T port map(A1 => n_293, A2 => n_1224, B1 => n_669, B2 => n_427, ZN => n_1099);
  g89704 : OAI22D0BWP7T port map(A1 => n_642, A2 => n_708, B1 => n_599, B2 => n_598, ZN => n_1170);
  g89702 : OAI22D0BWP7T port map(A1 => n_553, A2 => n_391, B1 => n_599, B2 => n_708, ZN => n_1135);
  g89449 : NR2D0BWP7T port map(A1 => n_688, A2 => n_597, ZN => n_834);
  g89448 : OAI221D0BWP7T port map(A1 => n_450, A2 => n_596, B1 => n_546, B2 => n_665, C => n_595, ZN => n_979);
  g89682 : MOAI22D0BWP7T port map(A1 => n_866, A2 => n_1052, B1 => n_1022, B2 => MISO_shift(41), ZN => n_594);
  g89502 : AOI221D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(12), B1 => n_681, B2 => n_225, C => n_404, ZN => n_593);
  g89503 : AO221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(49), B1 => n_1150, B2 => MISO_shift(48), C => n_469, Z => n_592);
  g89500 : OAI31D0BWP7T port map(A1 => n_496, A2 => n_985, A3 => n_667, B => n_233, ZN => n_591);
  g89675 : OAI22D0BWP7T port map(A1 => n_642, A2 => n_616, B1 => n_793, B2 => n_589, ZN => n_590);
  g89671 : MOAI22D0BWP7T port map(A1 => n_866, A2 => n_781, B1 => n_1150, B2 => MISO_shift(49), ZN => n_588);
  g89660 : INVD0BWP7T port map(I => n_586, ZN => n_587);
  g89550 : OAI22D0BWP7T port map(A1 => n_698, A2 => n_985, B1 => n_697, B2 => n_1117, ZN => n_585);
  g89536 : MOAI22D0BWP7T port map(A1 => n_583, A2 => n_1117, B1 => n_1022, B2 => MISO_shift(8), ZN => n_584);
  g89538 : MOAI22D0BWP7T port map(A1 => n_581, A2 => n_1052, B1 => n_876, B2 => n_1090, ZN => n_582);
  g89541 : OA32D1BWP7T port map(A1 => n_579, A2 => n_578, A3 => n_589, B1 => n_1013, B2 => n_581, Z => n_580);
  g89546 : MOAI22D0BWP7T port map(A1 => n_583, A2 => n_1010, B1 => n_1022, B2 => MISO_shift(5), ZN => n_577);
  g89547 : MOAI22D0BWP7T port map(A1 => n_697, A2 => n_1052, B1 => n_1022, B2 => MISO_shift(18), ZN => n_576);
  g89568 : OAI32D1BWP7T port map(A1 => n_901, A2 => n_567, A3 => n_575, B1 => n_604, B2 => n_638, ZN => n_938);
  g89570 : MOAI22D0BWP7T port map(A1 => n_572, A2 => n_637, B1 => n_574, B2 => n_551, ZN => n_1190);
  g89506 : OAI31D0BWP7T port map(A1 => MOSI_shift(2), A2 => n_464, A3 => n_506, B => n_461, ZN => n_1037);
  g89510 : OAI31D0BWP7T port map(A1 => n_465, A2 => n_365, A3 => n_771, B => n_481, ZN => n_728);
  g89511 : OAI32D1BWP7T port map(A1 => MOSI_shift(1), A2 => n_774, A3 => n_559, B1 => n_664, B2 => n_415, ZN => n_1032);
  g89522 : NR2D1BWP7T port map(A1 => n_395, A2 => n_467, ZN => n_1142);
  g89619 : OAI21D0BWP7T port map(A1 => n_497, A2 => n_538, B => n_646, ZN => n_878);
  g89614 : ND2D1BWP7T port map(A1 => n_573, A2 => n_572, ZN => n_898);
  g89532 : AOI21D0BWP7T port map(A1 => n_706, A2 => full_map_4_2(0), B => n_571, ZN => n_785);
  g89631 : OA21D0BWP7T port map(A1 => n_665, A2 => n_570, B => n_843, Z => n_822);
  g89696 : OAI22D0BWP7T port map(A1 => n_568, A2 => n_567, B1 => n_665, B2 => n_566, ZN => n_569);
  g89738 : INVD0BWP7T port map(I => n_564, ZN => n_565);
  g89740 : INVD0BWP7T port map(I => n_663, ZN => n_563);
  g89763 : NR2D0BWP7T port map(A1 => n_599, A2 => n_603, ZN => n_562);
  g89594 : AOI211XD0BWP7T port map(A1 => n_1022, A2 => MISO_shift(34), B => n_376, C => n_398, ZN => n_561);
  g89491 : AO222D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(72), B1 => n_352, B2 => n_272, C1 => n_1150, C2 => MISO_shift(71), Z => n_560);
  g89718 : MAOI22D0BWP7T port map(A1 => n_825, A2 => full_map_1_0(0), B1 => n_433, B2 => n_710, ZN => n_1096);
  g89720 : OAI22D0BWP7T port map(A1 => n_559, A2 => n_827, B1 => n_627, B2 => n_557, ZN => n_1024);
  g89721 : OAI22D0BWP7T port map(A1 => n_559, A2 => n_896, B1 => n_330, B2 => n_219, ZN => n_890);
  g89722 : MAOI22D0BWP7T port map(A1 => n_870, A2 => full_map_4_0(0), B1 => n_1231, B2 => n_558, ZN => n_712);
  g89725 : MOAI22D0BWP7T port map(A1 => n_665, A2 => n_557, B1 => n_556, B2 => n_514, ZN => n_926);
  g89700 : AOI22D0BWP7T port map(A1 => n_515, A2 => n_160, B1 => n_574, B2 => n_555, ZN => n_1073);
  g89519 : AOI222D0BWP7T port map(A1 => n_490, A2 => n_462, B1 => n_855, B2 => full_map_0_2(0), C1 => n_641, C2 => full_map_0_4(0), ZN => n_673);
  g89706 : MOAI22D0BWP7T port map(A1 => n_665, A2 => n_666, B1 => n_574, B2 => n_452, ZN => n_953);
  g89707 : MOAI22D0BWP7T port map(A1 => n_1231, A2 => n_554, B1 => n_870, B2 => full_map_5_14(0), ZN => n_626);
  g89712 : OAI22D0BWP7T port map(A1 => n_553, A2 => n_634, B1 => n_394, B2 => n_801, ZN => n_1169);
  g89516 : AOI31D0BWP7T port map(A1 => n_478, A2 => n_1086, A3 => full_map_12_14(0), B => n_406, ZN => n_1050);
  g89890 : OA21D0BWP7T port map(A1 => n_552, A2 => n_598, B => n_1215, Z => n_1163);
  g89713 : MAOI22D0BWP7T port map(A1 => n_870, A2 => full_map_5_0(0), B1 => n_1231, B2 => n_492, ZN => n_709);
  g89714 : AOI22D0BWP7T port map(A1 => n_869, A2 => n_551, B1 => n_870, B2 => full_map_3_14(0), ZN => n_586);
  g89733 : MOAI22D0BWP7T port map(A1 => n_1231, A2 => n_550, B1 => n_870, B2 => full_map_4_14(0), ZN => n_707);
  g89529 : NR2XD0BWP7T port map(A1 => n_723, A2 => n_511, ZN => n_738);
  g89777 : NR2XD0BWP7T port map(A1 => n_639, A2 => n_679, ZN => n_718);
  g89730 : MOAI22D0BWP7T port map(A1 => n_543, A2 => n_628, B1 => n_825, B2 => full_map_0_12(0), ZN => n_750);
  g89531 : IND2D1BWP7T port map(A1 => n_549, B1 => n_449, ZN => n_1091);
  g89895 : OAI21D0BWP7T port map(A1 => n_1224, A2 => n_548, B => n_547, ZN => n_769);
  g89734 : OA22D0BWP7T port map(A1 => n_456, A2 => n_487, B1 => n_546, B2 => n_545, Z => n_724);
  g89786 : NR2XD0BWP7T port map(A1 => n_853, A2 => n_679, ZN => n_787);
  g89683 : MOAI22D0BWP7T port map(A1 => n_543, A2 => n_567, B1 => n_542, B2 => full_map_0_12(0), ZN => n_544);
  g89537 : AOI22D0BWP7T port map(A1 => n_911, A2 => n_941, B1 => n_540, B2 => n_1086, ZN => n_541);
  g89542 : OAI32D0BWP7T port map(A1 => MOSI_shift(8), A2 => n_538, A3 => n_537, B1 => MOSI_shift(7), B2 => n_510, ZN => n_539);
  g89551 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(39), B1 => n_791, B2 => n_1009, ZN => n_536);
  g89555 : MOAI22D0BWP7T port map(A1 => n_595, A2 => n_1010, B1 => n_1022, B2 => MISO_shift(14), ZN => n_535);
  g89558 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(69), B1 => n_532, B2 => n_1009, ZN => n_534);
  g89561 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(54), B1 => n_532, B2 => n_833, ZN => n_533);
  g89562 : MAOI22D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(56), B1 => n_532, B2 => n_844, ZN => n_531);
  g89564 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(24), B1 => n_791, B2 => n_844, ZN => n_530);
  g89565 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(66), B1 => n_532, B2 => n_781, ZN => n_529);
  g89680 : AOI22D0BWP7T port map(A1 => n_556, A2 => full_map_1_0(0), B1 => n_635, B2 => full_map_1_14(0), ZN => n_528);
  g89668 : AO22D0BWP7T port map(A1 => n_825, A2 => n_675, B1 => n_526, B2 => n_641, Z => n_527);
  g89662 : AOI32D1BWP7T port map(A1 => n_524, A2 => n_523, A3 => full_map_0_11(0), B1 => n_825, B2 => full_map_0_13(0), ZN => n_525);
  g89584 : AOI31D0BWP7T port map(A1 => n_640, A2 => n_992, A3 => full_map_1_13(1), B => n_429, ZN => n_522);
  g89583 : INVD0BWP7T port map(I => n_721, ZN => n_521);
  g89581 : AOI32D1BWP7T port map(A1 => n_870, A2 => n_1087, A3 => full_map_0_13(0), B1 => n_520, B2 => n_519, ZN => n_998);
  g89578 : AOI32D1BWP7T port map(A1 => n_825, A2 => MOSI_shift(5), A3 => full_map_4_0(0), B1 => n_518, B2 => n_460, ZN => n_1000);
  g89576 : AOI33D1BWP7T port map(A1 => n_825, A2 => n_1017, A3 => full_map_4_14(0), B1 => n_870, B2 => n_1146, B3 => full_map_6_14(0), ZN => n_1144);
  g89602 : AOI32D1BWP7T port map(A1 => n_516, A2 => n_1090, A3 => full_map_5_0(0), B1 => n_517, B2 => full_map_3_0(0), ZN => n_1042);
  g89603 : AOI32D1BWP7T port map(A1 => n_516, A2 => n_1090, A3 => full_map_5_14(0), B1 => n_517, B2 => full_map_3_14(0), ZN => n_1184);
  g89609 : AOI31D0BWP7T port map(A1 => n_354, A2 => n_422, A3 => full_map_6_2(0), B => n_420, ZN => n_631);
  g89567 : AOI33D1BWP7T port map(A1 => n_515, A2 => n_514, A3 => n_513, B1 => n_542, B2 => n_1087, B3 => full_map_0_11(0), ZN => n_997);
  g89572 : AOI33D1BWP7T port map(A1 => n_869, A2 => n_512, A3 => n_67, B1 => n_870, B2 => n_637, B3 => full_map_2_0(0), ZN => n_1140);
  g89575 : AOI33D1BWP7T port map(A1 => n_804, A2 => n_524, A3 => full_map_0_9(0), B1 => n_825, B2 => n_1087, B3 => full_map_0_11(0), ZN => n_974);
  g89574 : AO33D0BWP7T port map(A1 => n_630, A2 => n_1080, A3 => full_map_14_11(0), B1 => n_804, B2 => n_353, B3 => full_map_0_5(0), Z => n_889);
  g89661 : INVD0BWP7T port map(I => n_736, ZN => n_782);
  g89615 : NR2D0BWP7T port map(A1 => n_511, A2 => n_619, ZN => n_763);
  g89534 : OAI21D0BWP7T port map(A1 => n_510, A2 => n_24, B => n_866, ZN => n_962);
  g89764 : NR2D0BWP7T port map(A1 => n_667, A2 => n_704, ZN => n_509);
  g89693 : AOI22D0BWP7T port map(A1 => n_760, A2 => n_941, B1 => n_1150, B2 => MISO_shift(24), ZN => n_508);
  g89694 : MOAI22D0BWP7T port map(A1 => n_506, A2 => n_662, B1 => n_505, B2 => full_map_14_10(0), ZN => n_507);
  g89697 : MOAI22D0BWP7T port map(A1 => n_729, A2 => n_446, B1 => n_706, B2 => full_map_0_3(0), ZN => n_504);
  g89870 : AOI22D0BWP7T port map(A1 => n_491, A2 => n_500, B1 => n_1150, B2 => MISO_shift(16), ZN => n_503);
  g89867 : AOI32D1BWP7T port map(A1 => n_239, A2 => n_158, A3 => full_map_1_13(1), B1 => n_501, B2 => n_500, ZN => n_502);
  g89864 : AOI22D0BWP7T port map(A1 => n_355, A2 => MOSI_shift(2), B1 => n_869, B2 => full_map_8_12(0), ZN => n_499);
  g89765 : NR2D0BWP7T port map(A1 => n_497, A2 => n_496, ZN => n_498);
  g89687 : MOAI22D0BWP7T port map(A1 => n_474, A2 => n_485, B1 => n_505, B2 => full_map_14_13(0), ZN => n_495);
  g89761 : ND2D0BWP7T port map(A1 => n_825, A2 => full_map_2_0(0), ZN => n_494);
  g89703 : AOI22D0BWP7T port map(A1 => n_520, A2 => n_1080, B1 => n_855, B2 => n_493, ZN => n_1159);
  g89724 : AOI22D0BWP7T port map(A1 => n_855, A2 => full_map_0_1(0), B1 => n_641, B2 => full_map_0_3(0), ZN => n_674);
  g89717 : AOI22D0BWP7T port map(A1 => n_515, A2 => n_454, B1 => n_855, B2 => full_map_0_0(0), ZN => n_1125);
  g89767 : ND2D0BWP7T port map(A1 => n_825, A2 => full_map_3_0(0), ZN => n_636);
  g89768 : ND2D1BWP7T port map(A1 => n_825, A2 => full_map_3_14(0), ZN => n_573);
  g89769 : NR2D0BWP7T port map(A1 => n_667, A2 => n_570, ZN => n_564);
  g89877 : AOI22D0BWP7T port map(A1 => n_869, A2 => n_159, B1 => n_453, B2 => n_916, ZN => n_1039);
  g89708 : MAOI22D0BWP7T port map(A1 => n_908, A2 => full_map_5_0(0), B1 => n_1224, B2 => n_492, ZN => n_625);
  g89710 : AOI22D0BWP7T port map(A1 => n_633, A2 => n_601, B1 => n_491, B2 => n_916, ZN => n_1083);
  g89711 : AO33D0BWP7T port map(A1 => n_869, A2 => n_512, A3 => n_519, B1 => n_490, B2 => n_489, B3 => n_967, Z => n_1055);
  g89772 : ND2D1BWP7T port map(A1 => n_870, A2 => full_map_1_14(0), ZN => n_646);
  g89728 : AOI22D0BWP7T port map(A1 => n_515, A2 => n_512, B1 => n_908, B2 => full_map_2_0(0), ZN => n_668);
  g89774 : NR2D0BWP7T port map(A1 => n_665, A2 => n_488, ZN => n_649);
  g89773 : NR2XD0BWP7T port map(A1 => n_497, A2 => n_488, ZN => n_655);
  g89737 : OAI22D0BWP7T port map(A1 => n_486, A2 => n_487, B1 => n_545, B2 => n_411, ZN => n_736);
  g89727 : MAOI22D0BWP7T port map(A1 => n_908, A2 => full_map_4_0(0), B1 => n_1224, B2 => n_418, ZN => n_671);
  g89732 : OAI22D0BWP7T port map(A1 => n_486, A2 => n_485, B1 => n_537, B2 => n_382, ZN => n_741);
  g89789 : NR2XD0BWP7T port map(A1 => n_667, A2 => n_965, ZN => n_663);
  g89794 : NR2XD0BWP7T port map(A1 => n_497, A2 => n_1052, ZN => n_660);
  g89735 : AOI22D0BWP7T port map(A1 => n_855, A2 => full_map_2_0(0), B1 => n_484, B2 => full_map_14_0(0), ZN => n_910);
  g89781 : ND2D1BWP7T port map(A1 => n_542, A2 => full_map_1_13(1), ZN => n_762);
  g89801 : ND2D1BWP7T port map(A1 => n_542, A2 => full_map_1_13(0), ZN => n_843);
  g89598 : ND2D1BWP7T port map(A1 => n_482, A2 => n_523, ZN => n_483);
  g89681 : AOI22D0BWP7T port map(A1 => n_484, A2 => full_map_14_2(0), B1 => n_480, B2 => full_map_14_4(0), ZN => n_481);
  g89679 : AOI22D0BWP7T port map(A1 => n_484, A2 => full_map_14_3(0), B1 => n_478, B2 => full_map_14_13(0), ZN => n_479);
  g89494 : OAI31D0BWP7T port map(A1 => n_1117, A2 => n_386, A3 => n_101, B => n_356, ZN => n_477);
  g89676 : AOI22D0BWP7T port map(A1 => n_706, A2 => n_60, B1 => n_1150, B2 => MISO_shift(47), ZN => n_476);
  g89504 : OAI221D0BWP7T port map(A1 => n_474, A2 => n_662, B1 => n_485, B2 => n_389, C => n_241, ZN => n_475);
  g89674 : AOI22D0BWP7T port map(A1 => n_855, A2 => n_526, B1 => n_1150, B2 => MISO_shift(18), ZN => n_473);
  g89673 : AOI22D0BWP7T port map(A1 => n_908, A2 => full_map_0_2(0), B1 => n_706, B2 => full_map_0_4(0), ZN => n_472);
  g89544 : AOI22D0BWP7T port map(A1 => n_706, A2 => n_526, B1 => n_540, B2 => n_941, ZN => n_471);
  g89672 : MAOI22D0BWP7T port map(A1 => n_484, A2 => full_map_14_4(0), B1 => n_405, B2 => n_432, ZN => n_470);
  g89669 : MOAI22D0BWP7T port map(A1 => n_435, A2 => n_468, B1 => n_876, B2 => n_1080, ZN => n_469);
  g89665 : OAI33D1BWP7T port map(A1 => n_466, A2 => n_1052, A3 => n_1224, B1 => n_465, B2 => n_464, B3 => n_1231, ZN => n_467);
  g89664 : AO32D1BWP7T port map(A1 => n_462, A2 => n_451, A3 => full_map_0_9(0), B1 => n_855, B2 => full_map_0_3(0), Z => n_463);
  g89663 : AOI32D0BWP7T port map(A1 => n_869, A2 => n_27, A3 => full_map_10_14(0), B1 => n_556, B2 => n_460, ZN => n_461);
  g89597 : NR2D0BWP7T port map(A1 => n_595, A2 => n_1052, ZN => n_459);
  g89517 : AOI31D0BWP7T port map(A1 => n_556, A2 => n_458, A3 => full_map_9_0(0), B => n_379, ZN => n_1063);
  g89883 : AOI22D0BWP7T port map(A1 => n_491, A2 => n_512, B1 => n_457, B2 => n_52, ZN => n_1043);
  g89604 : NR3D0BWP7T port map(A1 => n_456, A2 => MOSI_shift(2), A3 => n_596, ZN => n_571);
  g89605 : AOI31D0BWP7T port map(A1 => n_218, A2 => n_1146, A3 => full_map_4_0(0), B => n_371, ZN => n_779);
  g89608 : NR2XD0BWP7T port map(A1 => n_510, A2 => n_455, ZN => n_772);
  g89901 : INVD0BWP7T port map(I => n_866, ZN => n_715);
  MISO_shift_reg_3 : DFQD1BWP7T port map(CP => clk, D => n_372, Q => MISO_shift(3));
  MISO_shift_reg_12 : DFQD1BWP7T port map(CP => clk, D => n_359, Q => MISO_shift(12));
  g89880 : AOI22D0BWP7T port map(A1 => n_869, A2 => n_454, B1 => n_453, B2 => n_452, ZN => n_836);
  g89577 : AOI33D1BWP7T port map(A1 => n_855, A2 => n_967, A3 => full_map_0_4(0), B1 => n_337, B2 => n_451, B3 => full_map_14_10(0), ZN => n_690);
  g89573 : AOI32D1BWP7T port map(A1 => n_556, A2 => n_596, A3 => full_map_5_0(0), B1 => n_908, B2 => n_493, ZN => n_922);
  g89571 : OA33D0BWP7T port map(A1 => n_909, A2 => n_774, A3 => n_729, B1 => n_1010, B2 => n_388, B3 => n_771, Z => n_1115);
  MISO_shift_reg_9 : DFQD1BWP7T port map(CP => clk, D => n_358, Q => MISO_shift(9));
  g89600 : AOI21D0BWP7T port map(A1 => n_706, A2 => full_map_3_5(0), B => n_414, ZN => n_678);
  g89582 : OAI22D0BWP7T port map(A1 => n_450, A2 => n_417, B1 => n_605, B2 => n_546, ZN => n_688);
  g89632 : IOA21D1BWP7T port map(A1 => n_908, A2 => full_map_3_2(1), B => n_449, ZN => n_721);
  g89535 : OA221D0BWP7T port map(A1 => n_605, A2 => n_316, B1 => n_416, B2 => n_403, C => n_448, Z => n_933);
  g89685 : OAI22D0BWP7T port map(A1 => n_568, A2 => n_446, B1 => n_829, B2 => n_567, ZN => n_447);
  g89686 : MOAI22D0BWP7T port map(A1 => n_440, A2 => n_662, B1 => n_480, B2 => full_map_14_3(0), ZN => n_445);
  g89689 : MAOI22D0BWP7T port map(A1 => n_368, A2 => full_map_14_3(0), B1 => n_474, B2 => MOSI_shift(2), ZN => n_444);
  g89692 : AOI22D0BWP7T port map(A1 => n_795, A2 => n_820, B1 => n_1022, B2 => MISO_shift(43), ZN => n_443);
  g89684 : OAI22D0BWP7T port map(A1 => n_441, A2 => n_464, B1 => n_440, B2 => n_439, ZN => n_442);
  g89871 : MAOI22D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(19), B1 => n_552, B2 => n_437, ZN => n_438);
  g89868 : OAI22D0BWP7T port map(A1 => n_435, A2 => n_708, B1 => n_552, B2 => n_801, ZN => n_436);
  g89866 : OAI22D0BWP7T port map(A1 => n_771, A2 => n_708, B1 => n_433, B2 => n_432, ZN => n_434);
  g89865 : MAOI22D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(60), B1 => n_552, B2 => n_468, ZN => n_431);
  g89863 : MAOI22D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(25), B1 => n_448, B2 => n_1117, ZN => n_430);
  g89844 : OAI22D0BWP7T port map(A1 => n_428, A2 => n_427, B1 => n_435, B2 => n_437, ZN => n_429);
  g89846 : ND3D0BWP7T port map(A1 => n_501, A2 => n_596, A3 => full_map_7_10(0), ZN => n_426);
  g89849 : OAI31D0BWP7T port map(A1 => n_336, A2 => n_781, A3 => n_1224, B => n_235, ZN => n_425);
  g89850 : MOAI22D0BWP7T port map(A1 => n_428, A2 => n_468, B1 => n_1150, B2 => MISO_shift(45), ZN => n_424);
  g89851 : ND3D0BWP7T port map(A1 => n_491, A2 => n_422, A3 => full_map_1_13(0), ZN => n_423);
  g89857 : MAOI22D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(10), B1 => n_448, B2 => n_1013, ZN => n_421);
  g89861 : OAI22D0BWP7T port map(A1 => n_175, A2 => n_412, B1 => n_1231, B2 => n_11, ZN => n_420);
  g89874 : OAI22D0BWP7T port map(A1 => n_1224, A2 => n_419, B1 => n_1231, B2 => n_831, ZN => n_511);
  g89699 : OAI33D1BWP7T port map(A1 => n_418, A2 => n_1052, A3 => n_751, B1 => n_309, B2 => n_965, B3 => n_627, ZN => n_778);
  g89705 : OAI32D1BWP7T port map(A1 => n_301, A2 => n_417, A3 => n_537, B1 => n_416, B2 => n_387, ZN => n_549);
  g89766 : ND2D1BWP7T port map(A1 => n_855, A2 => full_map_3_0(0), ZN => n_572);
  g89715 : MOAI22D0BWP7T port map(A1 => n_575, A2 => n_628, B1 => n_641, B2 => full_map_0_2(0), ZN => n_602);
  g89716 : OAI33D1BWP7T port map(A1 => n_711, A2 => n_548, A3 => n_1224, B1 => n_566, B2 => n_893, B3 => n_415, ZN => n_952);
  g89723 : OAI22D0BWP7T port map(A1 => n_441, A2 => n_485, B1 => n_340, B2 => n_662, ZN => n_727);
  g89820 : CKND1BWP7T port map(I => n_414, ZN => n_583);
  g89729 : AO22D0BWP7T port map(A1 => n_396, A2 => n_629, B1 => MOSI_shift(2), B2 => n_413, Z => n_723);
  g89770 : ND2D1BWP7T port map(A1 => n_855, A2 => full_map_2_1(2), ZN => n_698);
  g89731 : AOI22D0BWP7T port map(A1 => n_480, A2 => full_map_11_4(0), B1 => n_413, B2 => n_367, ZN => n_765);
  g89736 : OAI22D0BWP7T port map(A1 => n_383, A2 => n_412, B1 => n_605, B2 => n_411, ZN => n_767);
  g89793 : ND2D1BWP7T port map(A1 => n_908, A2 => full_map_4_1(2), ZN => n_697);
  g89678 : MAOI22D0BWP7T port map(A1 => n_480, A2 => full_map_14_5(0), B1 => n_440, B2 => n_485, ZN => n_410);
  g89677 : MOAI22D0BWP7T port map(A1 => n_408, A2 => n_985, B1 => n_1150, B2 => MISO_shift(46), ZN => n_409);
  g89670 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(51), B1 => n_683, B2 => n_965, ZN => n_407);
  g89667 : OAI32D0BWP7T port map(A1 => n_263, A2 => n_1117, A3 => n_405, B1 => n_827, B2 => n_729, ZN => n_406);
  g89666 : MOAI22D0BWP7T port map(A1 => n_403, A2 => n_129, B1 => n_871, B2 => n_1015, ZN => n_404);
  g89589 : NR3D0BWP7T port map(A1 => n_486, A2 => n_401, A3 => MOSI_shift(2), ZN => n_402);
  g89900 : INVD0BWP7T port map(I => n_518, ZN => n_400);
  g89899 : INVD0BWP7T port map(I => n_398, ZN => n_399);
  g89587 : AOI32D1BWP7T port map(A1 => n_396, A2 => n_1015, A3 => n_31, B1 => n_1022, B2 => MISO_shift(67), ZN => n_397);
  g89585 : OAI32D0BWP7T port map(A1 => MOSI_shift(2), A2 => n_88, A3 => n_771, B1 => n_418, B2 => n_394, ZN => n_395);
  g89501 : OAI31D0BWP7T port map(A1 => n_679, A2 => n_901, A3 => n_405, B => n_329, ZN => n_393);
  g90018 : ND3D0BWP7T port map(A1 => n_869, A2 => n_40, A3 => full_map_10_11(0), ZN => n_392);
  g89885 : OAI22D0BWP7T port map(A1 => n_552, A2 => n_391, B1 => n_433, B2 => n_53, ZN => n_1114);
  g89879 : OAI22D0BWP7T port map(A1 => n_713, A2 => n_603, B1 => n_433, B2 => n_390, ZN => n_937);
  g89948 : CKND2D0BWP7T port map(A1 => n_869, A2 => n_916, ZN => n_547);
  g89569 : MAOI22D0BWP7T port map(A1 => n_295, A2 => n_749, B1 => n_389, B2 => n_89, ZN => n_607);
  g89881 : OAI32D1BWP7T port map(A1 => n_1010, A2 => n_708, A3 => n_339, B1 => n_672, B2 => n_748, ZN => n_692);
  g89886 : OAI22D0BWP7T port map(A1 => n_713, A2 => n_391, B1 => n_552, B2 => n_388, ZN => n_1046);
  MISO_shift_reg_6 : DFQD1BWP7T port map(CP => clk, D => n_349, Q => MISO_shift(6));
  g89891 : AOI32D1BWP7T port map(A1 => n_524, A2 => n_422, A3 => full_map_7_10(0), B1 => n_396, B2 => n_13, ZN => n_581);
  g89957 : ND2D0BWP7T port map(A1 => n_869, A2 => n_269, ZN => n_638);
  g89898 : MOAI22D0BWP7T port map(A1 => n_387, A2 => n_386, B1 => n_396, B2 => n_385, ZN => n_694);
  g89963 : ND2D1BWP7T port map(A1 => n_869, A2 => n_941, ZN => n_599);
  g89966 : ND2D1BWP7T port map(A1 => n_869, A2 => n_1086, ZN => n_669);
  g89905 : INVD1BWP7T port map(I => n_870, ZN => n_639);
  g89903 : INVD1BWP7T port map(I => n_635, ZN => n_642);
  g89906 : INVD1BWP7T port map(I => n_825, ZN => n_853);
  g89972 : ND2D1BWP7T port map(A1 => n_869, A2 => n_500, ZN => n_866);
  g89974 : ND2D1BWP7T port map(A1 => n_869, A2 => MOSI_shift(1), ZN => n_1215);
  g89869 : OAI22D0BWP7T port map(A1 => n_383, A2 => n_662, B1 => n_1224, B2 => n_382, ZN => n_384);
  g89759 : OAI21D0BWP7T port map(A1 => n_224, A2 => n_679, B => n_324, ZN => n_381);
  g89760 : NR2D0BWP7T port map(A1 => n_605, A2 => n_488, ZN => n_380);
  g89762 : INR2D0BWP7T port map(A1 => n_514, B1 => n_394, ZN => n_379);
  g89852 : MOAI22D0BWP7T port map(A1 => n_375, A2 => n_704, B1 => n_1150, B2 => MISO_shift(33), ZN => n_376);
  g89853 : MAOI22D0BWP7T port map(A1 => n_1150, A2 => MISO_shift(30), B1 => n_335, B2 => n_373, ZN => n_374);
  g89856 : AO221D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(3), B1 => n_1150, B2 => MISO_shift(2), C => n_286, Z => n_372);
  g89862 : OAI32D1BWP7T port map(A1 => n_37, A2 => n_965, A3 => n_751, B1 => n_664, B2 => n_627, ZN => n_371);
  g89739 : INVD0BWP7T port map(I => n_370, ZN => n_610);
  g89888 : IOA21D1BWP7T port map(A1 => n_524, A2 => full_map_0_13(0), B => n_568, ZN => n_482);
  g89889 : AOI22D0BWP7T port map(A1 => n_524, A2 => n_551, B1 => n_516, B2 => full_map_3_14(0), ZN => n_449);
  g89946 : NR2D0BWP7T port map(A1 => n_713, A2 => n_334, ZN => n_758);
  g89896 : MOAI22D0BWP7T port map(A1 => n_771, A2 => n_558, B1 => n_516, B2 => full_map_4_0(0), ZN => n_414);
  g89944 : NR2D0BWP7T port map(A1 => n_369, A2 => n_896, ZN => n_398);
  g89943 : NR2D0BWP7T port map(A1 => n_369, A2 => n_589, ZN => n_918);
  g89902 : INVD0BWP7T port map(I => n_556, ZN => n_553);
  g89882 : IOA21D1BWP7T port map(A1 => n_524, A2 => full_map_0_12(0), B => n_543, ZN => n_600);
  g89950 : NR2D1BWP7T port map(A1 => n_748, A2 => n_985, ZN => n_517);
  g89892 : MAOI22D0BWP7T port map(A1 => n_368, A2 => full_map_5_2(0), B1 => n_403, B2 => n_367, ZN => n_510);
  g89894 : OAI32D1BWP7T port map(A1 => n_546, A2 => n_416, A3 => n_578, B1 => n_412, B2 => n_273, ZN => n_911);
  full_map_reg_11_0_0 : DFQD1BWP7T port map(CP => clk, D => n_308, Q => full_map_11_0(0));
  full_map_reg_13_0_0 : DFQD1BWP7T port map(CP => clk, D => n_300, Q => full_map_13_0(0));
  full_map_reg_7_0_0 : DFQD1BWP7T port map(CP => clk, D => n_307, Q => full_map_7_0(0));
  g89951 : NR2XD0BWP7T port map(A1 => n_1231, A2 => n_366, ZN => n_518);
  g89785 : OR2D1BWP7T port map(A1 => n_545, A2 => n_496, Z => n_532);
  g89904 : INVD1BWP7T port map(I => n_706, ZN => n_497);
  g89897 : MAOI22D0BWP7T port map(A1 => n_516, A2 => full_map_4_14(0), B1 => n_771, B2 => n_550, ZN => n_595);
  g89975 : NR2XD0BWP7T port map(A1 => n_1231, A2 => n_833, ZN => n_635);
  g89961 : NR2D1BWP7T port map(A1 => n_1231, A2 => n_1009, ZN => n_574);
  g89962 : NR2D1BWP7T port map(A1 => n_1231, A2 => n_365, ZN => n_630);
  full_map_reg_14_2_0 : DFQD1BWP7T port map(CP => clk, D => n_319, Q => full_map_14_2(0));
  g89968 : NR2D1BWP7T port map(A1 => n_433, A2 => MOSI_shift(2), ZN => n_542);
  full_map_reg_8_0_0 : DFQD1BWP7T port map(CP => clk, D => n_321, Q => full_map_8_0(0));
  g89798 : IND2D1BWP7T port map(A1 => n_605, B1 => full_map_4_1(2), ZN => n_791);
  g89907 : INVD1BWP7T port map(I => n_855, ZN => n_667);
  full_map_reg_4_0_0 : DFQD1BWP7T port map(CP => clk, D => n_322, Q => full_map_4_0(0));
  g89908 : INVD1BWP7T port map(I => n_908, ZN => n_665);
  g89978 : NR2D1BWP7T port map(A1 => n_1231, A2 => n_455, ZN => n_870);
  g89979 : NR2D1BWP7T port map(A1 => n_1231, A2 => n_333, ZN => n_825);
  g89586 : AOI222D0BWP7T port map(A1 => n_363, A2 => n_1015, B1 => n_1150, B2 => MISO_shift(61), C1 => n_1022, C2 => MISO_shift(62), ZN => n_364);
  g89588 : ND4D0BWP7T port map(A1 => n_338, A2 => n_1090, A3 => MOSI_shift(2), A4 => MOSI_shift(7), ZN => n_362);
  g89591 : AOI222D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(71), B1 => n_360, B2 => n_1090, C1 => n_1150, C2 => MISO_shift(70), ZN => n_361);
  g89592 : OAI31D0BWP7T port map(A1 => n_1010, A2 => n_446, A3 => n_357, B => n_231, ZN => n_359);
  g89593 : OAI31D0BWP7T port map(A1 => n_985, A2 => n_628, A3 => n_357, B => n_230, ZN => n_358);
  g89595 : IND3D1BWP7T port map(A1 => n_545, B1 => full_map_5_6(0), B2 => n_820, ZN => n_356);
  g90046 : AOI21D0BWP7T port map(A1 => n_524, A2 => full_map_8_12(0), B => n_355, ZN => n_456);
  g90047 : AOI222D0BWP7T port map(A1 => n_524, A2 => full_map_0_10(0), B1 => n_354, B2 => full_map_0_2(0), C1 => n_353, C2 => full_map_0_6(0), ZN => n_559);
  full_map_reg_0_8_0 : DFQD1BWP7T port map(CP => clk, D => n_289, Q => full_map_0_8(0));
  full_map_reg_0_7_0 : DFQD1BWP7T port map(CP => clk, D => n_297, Q => full_map_0_7(0));
  full_map_reg_0_5_0 : DFQD1BWP7T port map(CP => clk, D => n_280, Q => full_map_0_5(0));
  full_map_reg_0_9_0 : DFQD1BWP7T port map(CP => clk, D => n_274, Q => full_map_0_9(0));
  full_map_reg_12_0_0 : DFQD1BWP7T port map(CP => clk, D => n_292, Q => full_map_12_0(0));
  full_map_reg_8_4_0 : DFQD1BWP7T port map(CP => clk, D => n_303, Q => full_map_8_4(0));
  full_map_reg_14_0_0 : DFQD1BWP7T port map(CP => clk, D => n_299, Q => full_map_14_0(0));
  full_map_reg_9_0_0 : DFQD1BWP7T port map(CP => clk, D => n_306, Q => full_map_9_0(0));
  full_map_reg_0_10_0 : DFQD1BWP7T port map(CP => clk, D => n_276, Q => full_map_0_10(0));
  full_map_reg_10_0_0 : DFQD1BWP7T port map(CP => clk, D => n_298, Q => full_map_10_0(0));
  full_map_reg_0_6_0 : DFQD1BWP7T port map(CP => clk, D => n_296, Q => full_map_0_6(0));
  full_map_reg_0_12_0 : DFQD1BWP7T port map(CP => clk, D => n_290, Q => full_map_0_12(0));
  full_map_reg_0_4_0 : DFQD1BWP7T port map(CP => clk, D => n_281, Q => full_map_0_4(0));
  full_map_reg_0_3_0 : DFQD1BWP7T port map(CP => clk, D => n_323, Q => full_map_0_3(0));
  full_map_reg_0_0_0 : DFQD1BWP7T port map(CP => clk, D => n_282, Q => full_map_0_0(0));
  full_map_reg_0_11_0 : DFQD1BWP7T port map(CP => clk, D => n_275, Q => full_map_0_11(0));
  full_map_reg_3_0_0 : DFQD1BWP7T port map(CP => clk, D => n_320, Q => full_map_3_0(0));
  full_map_reg_0_2_0 : DFQD1BWP7T port map(CP => clk, D => n_283, Q => full_map_0_2(0));
  full_map_reg_0_13_0 : DFQD1BWP7T port map(CP => clk, D => n_291, Q => full_map_0_13(0));
  full_map_reg_5_0_0 : DFQD1BWP7T port map(CP => clk, D => n_325, Q => full_map_5_0(0));
  full_map_reg_3_2_1 : DFQD1BWP7T port map(CP => clk, D => n_313, Q => full_map_3_2(1));
  g89989 : OAI31D0BWP7T port map(A1 => n_488, A2 => n_1013, A3 => n_567, B => n_226, ZN => n_352);
  g89982 : INVD0BWP7T port map(I => n_506, ZN => n_351);
  g89872 : AOI22D0BWP7T port map(A1 => n_363, A2 => n_941, B1 => n_1150, B2 => MISO_shift(64), ZN => n_350);
  g89859 : OAI21D0BWP7T port map(A1 => n_357, A2 => n_348, B => n_248, ZN => n_349);
  g89858 : AOI22D0BWP7T port map(A1 => n_360, A2 => n_1146, B1 => n_1022, B2 => MISO_shift(65), ZN => n_347);
  g89855 : AOI32D0BWP7T port map(A1 => n_515, A2 => n_820, A3 => n_345, B1 => n_1022, B2 => MISO_shift(26), ZN => n_346);
  g89854 : OAI32D1BWP7T port map(A1 => n_1, A2 => n_781, A3 => n_343, B1 => n_1010, B2 => n_383, ZN => n_344);
  g89845 : MOAI22D0BWP7T port map(A1 => n_270, A2 => n_86, B1 => n_1022, B2 => MISO_shift(1), ZN => n_342);
  g89771 : NR2XD0BWP7T port map(A1 => n_341, A2 => n_363, ZN => n_370);
  g89875 : MOAI22D0BWP7T port map(A1 => n_340, A2 => n_113, B1 => n_490, B2 => n_601, ZN => n_847);
  g89876 : AOI22D0BWP7T port map(A1 => n_368, A2 => full_map_8_4(0), B1 => n_240, B2 => full_map_8_12(0), ZN => n_450);
  g89887 : OAI33D1BWP7T port map(A1 => n_1009, A2 => n_34, A3 => n_339, B1 => n_465, B2 => n_111, B3 => n_343, ZN => n_377);
  g89942 : ND2D1BWP7T port map(A1 => n_338, A2 => n_385, ZN => n_857);
  g89726 : AOI33D1BWP7T port map(A1 => n_641, A2 => n_967, A3 => full_map_0_6(0), B1 => n_749, B2 => n_337, B3 => full_map_14_6(0), ZN => n_957);
  full_map_reg_11_14_0 : DFQD1BWP7T port map(CP => clk, D => n_221, Q => full_map_11_14(0));
  g89949 : NR2XD0BWP7T port map(A1 => n_1224, A2 => n_391, ZN => n_520);
  g89952 : NR2XD0BWP7T port map(A1 => n_537, A2 => n_336, ZN => n_619);
  g89953 : NR2D0BWP7T port map(A1 => n_335, A2 => n_567, ZN => n_1089);
  full_map_reg_8_14_0 : DFQD1BWP7T port map(CP => clk, D => n_249, Q => full_map_8_14(0));
  g89983 : INVD1BWP7T port map(I => n_575, ZN => n_633);
  g89893 : NR3D0BWP7T port map(A1 => n_335, A2 => n_367, A3 => MOSI_shift(8), ZN => n_540);
  g89958 : NR2D1BWP7T port map(A1 => n_335, A2 => n_446, ZN => n_876);
  g89965 : NR2D1BWP7T port map(A1 => n_1224, A2 => n_365, ZN => n_484);
  full_map_reg_4_14_0 : DFQD1BWP7T port map(CP => clk, D => n_260, Q => full_map_4_14(0));
  full_map_reg_7_10_0 : DFQD1BWP7T port map(CP => clk, D => n_257, Q => full_map_7_10(0));
  g89964 : NR2XD0BWP7T port map(A1 => n_335, A2 => n_334, ZN => n_760);
  g89973 : NR2XD0BWP7T port map(A1 => n_1224, A2 => n_833, ZN => n_556);
  g89977 : NR2XD0BWP7T port map(A1 => n_537, A2 => n_455, ZN => n_706);
  g89981 : NR2XD0BWP7T port map(A1 => n_1224, A2 => n_455, ZN => n_908);
  g89980 : NR2XD0BWP7T port map(A1 => n_1224, A2 => n_333, ZN => n_855);
  g90027 : IND3D0BWP7T port map(A1 => n_439, B1 => full_map_14_1(0), B2 => n_515, ZN => n_332);
  g90042 : AOI22D0BWP7T port map(A1 => n_524, A2 => full_map_14_9(0), B1 => n_353, B2 => full_map_14_5(0), ZN => n_330);
  g89590 : ND4D0BWP7T port map(A1 => n_368, A2 => n_1086, A3 => n_76, A4 => full_map_3_5(0), ZN => n_329);
  g90122 : INVD0BWP7T port map(I => n_435, ZN => n_328);
  g90020 : NR3D0BWP7T port map(A1 => n_1224, A2 => n_41, A3 => n_417, ZN => n_327);
  g90065 : INVD0BWP7T port map(I => n_552, ZN => n_453);
  g90064 : INVD1BWP7T port map(I => n_748, ZN => n_457);
  g90053 : AOI22D0BWP7T port map(A1 => n_271, A2 => full_map_10_8(0), B1 => n_524, B2 => full_map_10_12(0), ZN => n_486);
  g90123 : INVD1BWP7T port map(I => n_428, ZN => n_501);
  full_map_reg_7_14_0 : DFQD1BWP7T port map(CP => clk, D => n_259, Q => full_map_7_14(0));
  g90060 : INVD0BWP7T port map(I => n_326, ZN => n_505);
  full_map_reg_10_12_0 : DFQD1BWP7T port map(CP => clk, D => n_256, Q => full_map_10_12(0));
  full_map_reg_12_14_0 : DFQD1BWP7T port map(CP => clk, D => n_255, Q => full_map_12_14(0));
  g90124 : INVD0BWP7T port map(I => n_713, ZN => n_491);
  full_map_reg_9_14_0 : DFQD1BWP7T port map(CP => clk, D => n_258, Q => full_map_9_14(0));
  full_map_reg_6_14_0 : DFQD1BWP7T port map(CP => clk, D => n_265, Q => full_map_6_14(0));
  full_map_reg_10_14_0 : DFQD1BWP7T port map(CP => clk, D => n_262, Q => full_map_10_14(0));
  full_map_reg_13_14_0 : DFQD1BWP7T port map(CP => clk, D => n_254, Q => full_map_13_14(0));
  full_map_reg_5_14_0 : DFQD1BWP7T port map(CP => clk, D => n_238, Q => full_map_5_14(0));
  full_map_reg_10_11_0 : DFQD1BWP7T port map(CP => clk, D => n_266, Q => full_map_10_11(0));
  full_map_reg_3_5_0 : DFQD1BWP7T port map(CP => clk, D => n_247, Q => full_map_3_5(0));
  g90070 : INVD1BWP7T port map(I => n_1231, ZN => n_869);
  g89843 : ND2D0BWP7T port map(A1 => n_198, A2 => n_324, ZN => n_325);
  g89939 : ND2D0BWP7T port map(A1 => n_166, A2 => n_324, ZN => n_323);
  g89744 : ND2D0BWP7T port map(A1 => n_179, A2 => n_324, ZN => n_322);
  g89746 : ND2D0BWP7T port map(A1 => n_216, A2 => n_324, ZN => n_321);
  g89749 : ND2D0BWP7T port map(A1 => n_177, A2 => n_324, ZN => n_320);
  g89750 : ND2D0BWP7T port map(A1 => n_181, A2 => n_324, ZN => n_319);
  g89752 : OAI21D0BWP7T port map(A1 => n_131, A2 => n_411, B => n_324, ZN => n_318);
  g89754 : OAI21D0BWP7T port map(A1 => n_144, A2 => n_316, B => n_324, ZN => n_317);
  g89755 : OAI21D0BWP7T port map(A1 => n_155, A2 => n_579, B => n_324, ZN => n_315);
  g89756 : OAI21D0BWP7T port map(A1 => n_126, A2 => n_546, B => n_324, ZN => n_314);
  g89757 : ND2D0BWP7T port map(A1 => n_180, A2 => n_324, ZN => n_313);
  g89938 : OAI21D0BWP7T port map(A1 => n_152, A2 => n_570, B => n_324, ZN => n_312);
  g89821 : AOI222D0BWP7T port map(A1 => n_640, A2 => n_44, B1 => n_1150, B2 => MISO_shift(1), C1 => n_1022, C2 => MISO_shift(2), ZN => n_311);
  g89822 : OAI21D0BWP7T port map(A1 => n_125, A2 => n_309, B => n_324, ZN => n_310);
  g89823 : ND2D0BWP7T port map(A1 => n_211, A2 => n_324, ZN => n_308);
  g89824 : ND2D0BWP7T port map(A1 => n_209, A2 => n_324, ZN => n_307);
  g89826 : ND2D0BWP7T port map(A1 => n_205, A2 => n_324, ZN => n_306);
  g89936 : OAI21D0BWP7T port map(A1 => n_154, A2 => n_304, B => n_324, ZN => n_305);
  g89832 : ND2D0BWP7T port map(A1 => n_212, A2 => n_324, ZN => n_303);
  g89834 : OAI21D0BWP7T port map(A1 => n_121, A2 => n_301, B => n_324, ZN => n_302);
  g89836 : ND2D0BWP7T port map(A1 => n_196, A2 => n_324, ZN => n_300);
  g89838 : ND2D0BWP7T port map(A1 => n_184, A2 => n_324, ZN => n_299);
  g89842 : ND2D0BWP7T port map(A1 => n_183, A2 => n_324, ZN => n_298);
  g89935 : ND2D0BWP7T port map(A1 => n_200, A2 => n_324, ZN => n_297);
  g89933 : ND2D0BWP7T port map(A1 => n_167, A2 => n_324, ZN => n_296);
  g89847 : OAI21D0BWP7T port map(A1 => n_294, A2 => n_711, B => n_293, ZN => n_295);
  g89860 : ND2D0BWP7T port map(A1 => n_214, A2 => n_324, ZN => n_292);
  g89932 : ND2D0BWP7T port map(A1 => n_203, A2 => n_324, ZN => n_291);
  g89909 : ND2D0BWP7T port map(A1 => n_210, A2 => n_324, ZN => n_290);
  g89910 : ND2D0BWP7T port map(A1 => n_161, A2 => n_324, ZN => n_289);
  g89911 : OAI21D0BWP7T port map(A1 => n_122, A2 => n_287, B => n_324, ZN => n_288);
  g89912 : INR2D0BWP7T port map(A1 => n_285, B1 => n_357, ZN => n_286);
  g89914 : OAI21D0BWP7T port map(A1 => n_123, A2 => n_566, B => n_324, ZN => n_284);
  g89915 : ND2D0BWP7T port map(A1 => n_172, A2 => n_324, ZN => n_283);
  g89919 : ND2D0BWP7T port map(A1 => n_201, A2 => n_324, ZN => n_282);
  g89921 : ND2D0BWP7T port map(A1 => n_168, A2 => n_324, ZN => n_281);
  g89925 : ND2D0BWP7T port map(A1 => n_170, A2 => n_324, ZN => n_280);
  g89878 : OAI22D0BWP7T port map(A1 => n_829, A2 => n_279, B1 => n_751, B2 => MOSI_shift(1), ZN => n_608);
  g89947 : ND2D0BWP7T port map(A1 => n_641, A2 => full_map_3_2(1), ZN => n_408);
  g89940 : NR2D0BWP7T port map(A1 => n_387, A2 => MOSI_shift(7), ZN => n_413);
  g89954 : ND2D0BWP7T port map(A1 => n_515, A2 => n_941, ZN => n_394);
  full_map_reg_14_8_0 : DFQD1BWP7T port map(CP => clk, D => n_215, Q => full_map_14_8(0));
  full_map_reg_14_6_0 : DFQD1BWP7T port map(CP => clk, D => n_185, Q => full_map_14_6(0));
  full_map_reg_14_11_0 : DFQD1BWP7T port map(CP => clk, D => n_190, Q => full_map_14_11(0));
  g90030 : OAI21D0BWP7T port map(A1 => n_223, A2 => n_222, B => n_324, ZN => n_278);
  g90021 : MAOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(11), B1 => n_405, B2 => n_621, ZN => n_277);
  g89986 : ND2D0BWP7T port map(A1 => n_164, A2 => n_324, ZN => n_276);
  g89984 : ND2D0BWP7T port map(A1 => n_165, A2 => n_324, ZN => n_275);
  g89985 : ND2D0BWP7T port map(A1 => n_162, A2 => n_324, ZN => n_274);
  g90098 : ND2D1BWP7T port map(A1 => n_524, A2 => n_629, ZN => n_326);
  g90058 : INVD0BWP7T port map(I => n_273, ZN => n_355);
  g90049 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_0_4(0), B1 => n_271, B2 => full_map_0_8(0), ZN => n_543);
  g90050 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_14_5(0), B1 => n_271, B2 => full_map_14_9(0), ZN => n_474);
  g90051 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_14_7(0), B1 => n_271, B2 => full_map_14_11(0), ZN => n_440);
  g90052 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_14_4(0), B1 => n_271, B2 => full_map_14_8(0), ZN => n_506);
  g89956 : NR2XD0BWP7T port map(A1 => n_270, A2 => n_662, ZN => n_795);
  g90063 : INVD0BWP7T port map(I => n_335, ZN => n_681);
  g89955 : ND2D1BWP7T port map(A1 => n_641, A2 => full_map_2_1(2), ZN => n_683);
  g90095 : ND2D1BWP7T port map(A1 => n_524, A2 => full_map_1_13(0), ZN => n_369);
  g90096 : ND2D1BWP7T port map(A1 => n_524, A2 => full_map_1_13(1), ZN => n_904);
  full_map_reg_14_7_0 : DFQD1BWP7T port map(CP => clk, D => n_186, Q => full_map_14_7(0));
  g90048 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_14_6(0), B1 => n_271, B2 => full_map_14_10(0), ZN => n_441);
  g90055 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_0_6(0), B1 => n_271, B2 => full_map_0_10(0), ZN => n_575);
  g89960 : ND2D0BWP7T port map(A1 => n_515, A2 => n_269, ZN => n_802);
  full_map_reg_5_6_0 : DFQD1BWP7T port map(CP => clk, D => n_204, Q => full_map_5_6(0));
  g90054 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_0_5(0), B1 => n_271, B2 => full_map_0_9(0), ZN => n_568);
  g90097 : ND2D1BWP7T port map(A1 => n_524, A2 => n_500, ZN => n_448);
  full_map_reg_14_10_0 : DFQD1BWP7T port map(CP => clk, D => n_193, Q => full_map_14_10(0));
  g90100 : NR2XD0BWP7T port map(A1 => n_195, A2 => n_301, ZN => n_396);
  full_map_reg_14_4_0 : DFQD1BWP7T port map(CP => clk, D => n_192, Q => full_map_14_4(0));
  full_map_reg_10_8_0 : DFQD1BWP7T port map(CP => clk, D => n_189, Q => full_map_10_8(0));
  full_map_reg_14_5_0 : DFQD1BWP7T port map(CP => clk, D => n_191, Q => full_map_14_5(0));
  full_map_reg_14_9_0 : DFQD1BWP7T port map(CP => clk, D => n_207, Q => full_map_14_9(0));
  g90172 : ND2D1BWP7T port map(A1 => n_524, A2 => n_941, ZN => n_435);
  g90174 : ND2D1BWP7T port map(A1 => n_524, A2 => n_1015, ZN => n_428);
  bit_counter_reg_1 : DFQD1BWP7T port map(CP => clk, D => n_173, Q => bit_counter(1));
  full_map_reg_6_0_0 : DFKSND1BWP7T port map(CP => clk, D => n_5, SN => n_145, Q => UNCONNECTED, QN => full_map_6_0(0));
  g89967 : NR2D1BWP7T port map(A1 => n_270, A2 => n_412, ZN => n_871);
  full_map_reg_14_3_0 : DFQD1BWP7T port map(CP => clk, D => n_187, Q => full_map_14_3(0));
  g89969 : ND2D1BWP7T port map(A1 => n_368, A2 => n_268, ZN => n_545);
  g90066 : CKND1BWP7T port map(I => n_516, ZN => n_433);
  g90056 : AOI22D0BWP7T port map(A1 => n_272, A2 => full_map_0_7(0), B1 => n_271, B2 => full_map_0_11(0), ZN => n_729);
  g90175 : ND2D1BWP7T port map(A1 => n_524, A2 => n_1086, ZN => n_713);
  g89971 : ND2D1BWP7T port map(A1 => n_515, A2 => n_268, ZN => n_605);
  g90109 : ND2D1BWP7T port map(A1 => n_524, A2 => n_820, ZN => n_552);
  g90108 : ND2D1BWP7T port map(A1 => n_524, A2 => n_38, ZN => n_748);
  g89976 : ND2D1BWP7T port map(A1 => n_515, A2 => n_909, ZN => n_1239);
  g90121 : ND2D1BWP7T port map(A1 => n_524, A2 => MOSI_shift(2), ZN => n_1231);
  g90025 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(27), B1 => n_1150, B2 => MISO_shift(26), ZN => n_267);
  g89743 : ND2D0BWP7T port map(A1 => n_151, A2 => n_324, ZN => n_266);
  g89745 : ND2D0BWP7T port map(A1 => n_136, A2 => n_324, ZN => n_265);
  g89747 : OAI21D0BWP7T port map(A1 => n_94, A2 => n_263, B => n_324, ZN => n_264);
  g89748 : ND2D0BWP7T port map(A1 => n_134, A2 => n_324, ZN => n_262);
  g89751 : OAI21D0BWP7T port map(A1 => n_95, A2 => n_432, B => n_324, ZN => n_261);
  g89753 : ND2D0BWP7T port map(A1 => n_138, A2 => n_324, ZN => n_260);
  g89827 : ND2D0BWP7T port map(A1 => n_140, A2 => n_324, ZN => n_259);
  g89828 : ND2D0BWP7T port map(A1 => n_141, A2 => n_324, ZN => n_258);
  g89831 : ND2D0BWP7T port map(A1 => n_150, A2 => n_324, ZN => n_257);
  g89833 : ND2D0BWP7T port map(A1 => n_147, A2 => n_324, ZN => n_256);
  g89835 : ND2D0BWP7T port map(A1 => n_157, A2 => n_324, ZN => n_255);
  g89837 : ND2D0BWP7T port map(A1 => n_146, A2 => n_324, ZN => n_254);
  g89839 : OAI21D0BWP7T port map(A1 => n_91, A2 => n_252, B => n_324, ZN => n_253);
  g89840 : OAI21D0BWP7T port map(A1 => n_115, A2 => n_465, B => n_324, ZN => n_251);
  g89841 : ND2D0BWP7T port map(A1 => n_149, A2 => n_324, ZN => n_250);
  g89742 : ND2D0BWP7T port map(A1 => n_137, A2 => n_324, ZN => n_249);
  g90024 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(6), B1 => n_1150, B2 => MISO_shift(5), ZN => n_248);
  g89922 : ND2D0BWP7T port map(A1 => n_130, A2 => n_324, ZN => n_247);
  g89926 : OAI21D0BWP7T port map(A1 => n_75, A2 => n_538, B => n_324, ZN => n_246);
  g89929 : OAI21D0BWP7T port map(A1 => n_96, A2 => n_244, B => n_324, ZN => n_245);
  g90010 : NR3D0BWP7T port map(A1 => n_771, A2 => n_1117, A3 => n_492, ZN => n_243);
  g89987 : AO211D0BWP7T port map(A1 => n_58, A2 => bit_counter(2), B => n_102, C => n_99, Z => n_242);
  g89996 : ND3D0BWP7T port map(A1 => n_749, A2 => n_458, A3 => full_map_14_1(0), ZN => n_241);
  g89884 : AO33D0BWP7T port map(A1 => n_240, A2 => n_551, A3 => n_1090, B1 => n_239, B2 => n_451, B3 => full_map_0_10(0), Z => n_691);
  g89941 : NR2D0BWP7T port map(A1 => n_127, A2 => n_416, ZN => n_341);
  g90082 : NR2D0BWP7T port map(A1 => n_771, A2 => n_427, ZN => n_597);
  g89873 : AOI33D1BWP7T port map(A1 => n_240, A2 => n_35, A3 => n_1086, B1 => n_478, B2 => n_820, B3 => full_map_13_14(0), ZN => n_846);
  g89830 : ND2D0BWP7T port map(A1 => n_143, A2 => n_324, ZN => n_238);
  g90034 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(38), B1 => n_1150, B2 => MISO_shift(37), ZN => n_237);
  g90035 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(56), B1 => n_1150, B2 => MISO_shift(55), ZN => n_236);
  g90036 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(23), B1 => n_1150, B2 => MISO_shift(22), ZN => n_235);
  g90037 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(60), B1 => n_1150, B2 => MISO_shift(59), ZN => n_234);
  g90038 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(30), B1 => n_1150, B2 => MISO_shift(29), ZN => n_233);
  g90039 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(33), B1 => n_1150, B2 => MISO_shift(32), ZN => n_232);
  g90040 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(12), B1 => n_1150, B2 => MISO_shift(11), ZN => n_231);
  g90041 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(9), B1 => n_1150, B2 => MISO_shift(8), ZN => n_230);
  g90043 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(32), B1 => n_1150, B2 => MISO_shift(31), ZN => n_229);
  g90032 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(15), B1 => n_1150, B2 => MISO_shift(14), ZN => n_228);
  g90029 : AOI22D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(40), B1 => n_1150, B2 => MISO_shift(39), ZN => n_227);
  g90161 : AOI32D0BWP7T port map(A1 => n_422, A2 => n_1015, A3 => full_map_4_1(2), B1 => n_225, B2 => full_map_1_1(2), ZN => n_226);
  g90079 : CKAN2D0BWP7T port map(A1 => n_223, A2 => n_222, Z => n_224);
  g89825 : ND2D0BWP7T port map(A1 => n_117, A2 => n_324, ZN => n_221);
  g90129 : MAOI22D0BWP7T port map(A1 => n_804, A2 => full_map_0_1(0), B1 => n_219, B2 => n_2, ZN => n_220);
  MOSI_shift_reg_0 : DFQD1BWP7T port map(CP => clk, D => n_153, Q => MOSI_shift(0));
  g90057 : INVD1BWP7T port map(I => n_218, ZN => n_415);
  g90092 : ND2D1BWP7T port map(A1 => n_272, A2 => full_map_8_4(0), ZN => n_273);
  g90068 : INVD0BWP7T port map(I => n_641, ZN => n_375);
  g90061 : INVD0BWP7T port map(I => n_270, ZN => n_338);
  g90094 : ND2D1BWP7T port map(A1 => n_272, A2 => full_map_5_6(0), ZN => n_403);
  g90062 : INVD1BWP7T port map(I => n_217, ZN => n_627);
  g90107 : ND2D1BWP7T port map(A1 => n_272, A2 => full_map_3_5(0), ZN => n_335);
  g90067 : INVD1BWP7T port map(I => n_368, ZN => n_537);
  g90110 : NR2D1BWP7T port map(A1 => n_771, A2 => n_455, ZN => n_516);
  state_reg_0 : DFQD1BWP7T port map(CP => clk, D => n_156, Q => state(0));
  g90069 : INVD1BWP7T port map(I => n_515, ZN => n_1224);
  g90015 : OAI21D0BWP7T port map(A1 => n_213, A2 => n_487, B => full_map_8_0(0), ZN => n_216);
  g89924 : ND2D0BWP7T port map(A1 => n_110, A2 => n_324, ZN => n_215);
  g90011 : OAI21D0BWP7T port map(A1 => n_213, A2 => n_485, B => full_map_12_0(0), ZN => n_214);
  g89992 : OAI21D0BWP7T port map(A1 => n_1259, A2 => n_833, B => full_map_8_4(0), ZN => n_212);
  g90009 : OAI21D0BWP7T port map(A1 => n_208, A2 => n_487, B => full_map_11_0(0), ZN => n_211);
  g90157 : OAI21D0BWP7T port map(A1 => n_827, A2 => n_202, B => full_map_0_12(0), ZN => n_210);
  g90008 : OAI21D0BWP7T port map(A1 => n_208, A2 => n_416, B => full_map_7_0(0), ZN => n_209);
  g89913 : ND2D0BWP7T port map(A1 => n_103, A2 => n_324, ZN => n_207);
  g89741 : ND2D0BWP7T port map(A1 => n_97, A2 => n_324, ZN => n_206);
  g90006 : OAI21D0BWP7T port map(A1 => n_197, A2 => n_487, B => full_map_9_0(0), ZN => n_205);
  g89758 : ND2D0BWP7T port map(A1 => n_98, A2 => n_324, ZN => n_204);
  g90153 : OAI21D0BWP7T port map(A1 => n_896, A2 => n_202, B => full_map_0_13(0), ZN => n_203);
  g90143 : OAI21D0BWP7T port map(A1 => n_827, A2 => n_171, B => full_map_0_0(0), ZN => n_201);
  g90150 : OAI21D0BWP7T port map(A1 => n_348, A2 => n_169, B => full_map_0_7(0), ZN => n_200);
  g89829 : OAI21D0BWP7T port map(A1 => n_62, A2 => n_496, B => n_324, ZN => n_199);
  g90004 : OAI21D0BWP7T port map(A1 => n_197, A2 => n_416, B => full_map_5_0(0), ZN => n_198);
  g90001 : OAI21D0BWP7T port map(A1 => n_197, A2 => n_485, B => full_map_13_0(0), ZN => n_196);
  g90179 : INVD0BWP7T port map(I => n_272, ZN => n_195);
  g89916 : ND2D0BWP7T port map(A1 => n_114, A2 => n_324, ZN => n_194);
  g89918 : ND2D0BWP7T port map(A1 => n_90, A2 => n_324, ZN => n_193);
  g89920 : ND2D0BWP7T port map(A1 => n_83, A2 => n_324, ZN => n_192);
  g89923 : ND2D0BWP7T port map(A1 => n_80, A2 => n_324, ZN => n_191);
  g89927 : ND2D0BWP7T port map(A1 => n_92, A2 => n_324, ZN => n_190);
  g89928 : ND2D0BWP7T port map(A1 => n_87, A2 => n_324, ZN => n_189);
  g89930 : ND2D0BWP7T port map(A1 => n_108, A2 => n_324, ZN => n_188);
  g89931 : ND2D0BWP7T port map(A1 => n_112, A2 => n_324, ZN => n_187);
  g89934 : ND2D0BWP7T port map(A1 => n_82, A2 => n_324, ZN => n_186);
  g89937 : ND2D0BWP7T port map(A1 => n_81, A2 => n_324, ZN => n_185);
  g89997 : OAI21D0BWP7T port map(A1 => n_182, A2 => n_485, B => full_map_14_0(0), ZN => n_184);
  g89999 : OAI21D0BWP7T port map(A1 => n_182, A2 => n_487, B => full_map_10_0(0), ZN => n_183);
  MOSI_shift_reg_9 : DFQD1BWP7T port map(CP => clk, D => n_72, Q => MOSI_shift(9));
  g90102 : NR2D1BWP7T port map(A1 => n_751, A2 => n_391, ZN => n_363);
  g90099 : ND2D1BWP7T port map(A1 => n_271, A2 => full_map_1_13(0), ZN => n_357);
  g90114 : NR2D1BWP7T port map(A1 => n_751, A2 => n_628, ZN => n_641);
  g90181 : INVD1BWP7T port map(I => n_771, ZN => n_524);
  g90019 : OAI21D0BWP7T port map(A1 => n_182, A2 => n_662, B => full_map_14_2(0), ZN => n_181);
  g90022 : OAI21D0BWP7T port map(A1 => n_208, A2 => n_446, B => full_map_3_2(1), ZN => n_180);
  g90026 : OAI21D0BWP7T port map(A1 => n_213, A2 => n_416, B => full_map_4_0(0), ZN => n_179);
  g90160 : AO21D0BWP7T port map(A1 => n_104, A2 => bit_counter(0), B => n_71, Z => n_178);
  g90017 : OAI21D0BWP7T port map(A1 => n_208, A2 => n_567, B => full_map_3_0(0), ZN => n_177);
  g90080 : ND2D0BWP7T port map(A1 => n_1022, A2 => MISO_shift(48), ZN => n_176);
  g90088 : CKND2D0BWP7T port map(A1 => n_271, A2 => full_map_10_8(0), ZN => n_175);
  g90081 : NR2D0BWP7T port map(A1 => n_632, A2 => n_546, ZN => n_174);
  g90158 : OAI31D0BWP7T port map(A1 => bit_counter(1), A2 => n_7, A3 => n_106, B => n_100, ZN => n_173);
  g90151 : OAI21D0BWP7T port map(A1 => n_279, A2 => n_171, B => full_map_0_2(0), ZN => n_172);
  g90149 : OAI21D0BWP7T port map(A1 => n_896, A2 => n_169, B => full_map_0_5(0), ZN => n_170);
  g90144 : OAI21D0BWP7T port map(A1 => n_827, A2 => n_169, B => full_map_0_4(0), ZN => n_168);
  g90142 : OAI21D0BWP7T port map(A1 => n_279, A2 => n_169, B => full_map_0_6(0), ZN => n_167);
  g90139 : OAI21D0BWP7T port map(A1 => n_348, A2 => n_171, B => full_map_0_3(0), ZN => n_166);
  g90131 : OAI21D0BWP7T port map(A1 => n_348, A2 => n_1260, B => full_map_0_11(0), ZN => n_165);
  g90133 : OAI21D0BWP7T port map(A1 => n_279, A2 => n_1260, B => full_map_0_10(0), ZN => n_164);
  g90134 : OAI21D0BWP7T port map(A1 => n_896, A2 => n_1260, B => full_map_0_9(0), ZN => n_162);
  g90137 : OAI21D0BWP7T port map(A1 => n_827, A2 => n_1260, B => full_map_0_8(0), ZN => n_161);
  g90044 : AOI21D0BWP7T port map(A1 => n_512, A2 => n_269, B => n_160, ZN => n_730);
  g90105 : NR2XD0BWP7T port map(A1 => n_751, A2 => n_333, ZN => n_217);
  g90045 : IAO21D0BWP7T port map(A1 => n_548, A2 => n_366, B => n_159, ZN => n_293);
  g90089 : NR2XD0BWP7T port map(A1 => n_751, A2 => n_455, ZN => n_218);
  g90166 : AOI22D0BWP7T port map(A1 => n_158, A2 => full_map_14_12(0), B1 => n_451, B2 => full_map_14_8(0), ZN => n_340);
  g90170 : AOI22D0BWP7T port map(A1 => n_158, A2 => full_map_10_12(0), B1 => n_451, B2 => full_map_10_8(0), ZN => n_383);
  g90171 : AO22D0BWP7T port map(A1 => n_158, A2 => full_map_0_12(0), B1 => full_map_0_8(0), B2 => n_451, Z => n_490);
  g90091 : ND2D1BWP7T port map(A1 => n_271, A2 => full_map_7_10(0), ZN => n_387);
  g90093 : INR2D0BWP7T port map(A1 => full_map_3_2(1), B1 => n_632, ZN => n_360);
  g90103 : ND2D1BWP7T port map(A1 => n_271, A2 => full_map_10_11(0), ZN => n_270);
  g90104 : NR2D1BWP7T port map(A1 => n_751, A2 => n_662, ZN => n_480);
  g90111 : NR2XD0BWP7T port map(A1 => n_751, A2 => n_367, ZN => n_368);
  MOSI_shift_reg_4 : DFQD1BWP7T port map(CP => clk, D => n_107, Q => MOSI_shift(4));
  g90120 : NR2D1BWP7T port map(A1 => n_751, A2 => MOSI_shift(2), ZN => n_515);
  g90000 : OAI21D0BWP7T port map(A1 => n_148, A2 => n_662, B => full_map_12_14(0), ZN => n_157);
  g89596 : OAI21D0BWP7T port map(A1 => n_49, A2 => reset, B => n_23, ZN => n_156);
  g90074 : NR2XD0BWP7T port map(A1 => n_182, A2 => n_446, ZN => n_155);
  g90185 : NR2D0BWP7T port map(A1 => n_279, A2 => n_202, ZN => n_154);
  g89848 : AO32D1BWP7T port map(A1 => n_50, A2 => n_66, A3 => MOSI, B1 => n_51, B2 => MOSI_shift(0), Z => n_153);
  g90221 : NR2D0BWP7T port map(A1 => n_373, A2 => n_171, ZN => n_152);
  g89990 : OAI31D0BWP7T port map(A1 => n_412, A2 => n_1010, A3 => n_1260, B => full_map_10_11(0), ZN => n_151);
  g89991 : OAI31D0BWP7T port map(A1 => n_1052, A2 => n_386, A3 => n_1260, B => full_map_7_10(0), ZN => n_150);
  g89993 : OAI21D0BWP7T port map(A1 => n_148, A2 => n_487, B => full_map_8_12(0), ZN => n_149);
  g89994 : OAI21D0BWP7T port map(A1 => n_135, A2 => n_487, B => full_map_10_12(0), ZN => n_147);
  g89995 : OAI21D0BWP7T port map(A1 => n_142, A2 => n_662, B => full_map_13_14(0), ZN => n_146);
  g89998 : AO21D0BWP7T port map(A1 => n_54, A2 => n_422, B => full_map_6_0(0), Z => n_145);
  g90071 : NR2D0BWP7T port map(A1 => n_197, A2 => n_386, ZN => n_144);
  g90002 : OAI21D0BWP7T port map(A1 => n_142, A2 => n_386, B => full_map_5_14(0), ZN => n_143);
  g90003 : OAI21D0BWP7T port map(A1 => n_142, A2 => n_412, B => full_map_9_14(0), ZN => n_141);
  g90005 : OAI21D0BWP7T port map(A1 => n_116, A2 => n_386, B => full_map_7_14(0), ZN => n_140);
  g90176 : INVD0BWP7T port map(I => n_640, ZN => n_139);
  g90012 : OAI21D0BWP7T port map(A1 => n_148, A2 => n_386, B => full_map_4_14(0), ZN => n_138);
  g90013 : OAI21D0BWP7T port map(A1 => n_148, A2 => n_412, B => full_map_8_14(0), ZN => n_137);
  g90014 : OAI21D0BWP7T port map(A1 => n_135, A2 => n_386, B => full_map_6_14(0), ZN => n_136);
  g90016 : OAI21D0BWP7T port map(A1 => n_135, A2 => n_412, B => full_map_10_14(0), ZN => n_134);
  g90023 : ND4D0BWP7T port map(A1 => n_353, A2 => n_85, A3 => n_1146, A4 => full_map_3_5(0), ZN => n_133);
  g90031 : ND4D0BWP7T port map(A1 => n_354, A2 => n_1015, A3 => n_345, A4 => n_367, ZN => n_132);
  MOSI_shift_reg_12 : DFQD1BWP7T port map(CP => clk, D => n_56, Q => MOSI_shift(12));
  g90173 : AOI22D0BWP7T port map(A1 => n_354, A2 => full_map_0_3(0), B1 => n_353, B2 => full_map_0_7(0), ZN => n_829);
  g90126 : NR2XD0BWP7T port map(A1 => n_182, A2 => n_386, ZN => n_131);
  g90146 : OAI21D0BWP7T port map(A1 => n_129, A2 => n_169, B => full_map_3_5(0), ZN => n_130);
  g90127 : OAI22D0BWP7T port map(A1 => n_548, A2 => n_844, B1 => n_419, B2 => n_833, ZN => n_128);
  g90162 : AOI22D0BWP7T port map(A1 => n_354, A2 => full_map_5_2(0), B1 => n_353, B2 => full_map_5_6(0), ZN => n_127);
  g90072 : NR2XD0BWP7T port map(A1 => n_213, A2 => n_386, ZN => n_126);
  g90128 : NR2XD0BWP7T port map(A1 => n_182, A2 => n_567, ZN => n_125);
  g90163 : AO22D0BWP7T port map(A1 => n_354, A2 => full_map_14_2(0), B1 => full_map_14_6(0), B2 => n_353, Z => n_124);
  g90210 : NR2D0BWP7T port map(A1 => n_896, A2 => n_171, ZN => n_123);
  g90211 : NR2D0BWP7T port map(A1 => n_589, A2 => n_171, ZN => n_122);
  g90078 : NR2XD0BWP7T port map(A1 => n_1259, A2 => n_1052, ZN => n_121);
  g90125 : MOAI22D0BWP7T port map(A1 => n_548, A2 => n_833, B1 => n_118, B2 => n_1146, ZN => n_119);
  g90007 : OAI21D0BWP7T port map(A1 => n_116, A2 => n_412, B => full_map_11_14(0), ZN => n_117);
  MOSI_shift_reg_13 : DFQD1BWP7T port map(CP => clk, D => n_61, Q => MOSI_shift(13));
  MOSI_shift_reg_10 : DFQD1BWP7T port map(CP => clk, D => n_59, Q => MOSI_shift(10));
  MOSI_shift_reg_11 : DFQD1BWP7T port map(CP => clk, D => n_65, Q => MOSI_shift(11));
  g90165 : AOI22D0BWP7T port map(A1 => n_354, A2 => full_map_14_3(0), B1 => n_353, B2 => full_map_14_7(0), ZN => n_389);
  g90188 : NR2XD0BWP7T port map(A1 => n_373, A2 => n_202, ZN => n_223);
  g90177 : CKND0BWP7T port map(I => n_240, ZN => n_339);
  bit_counter_reg_3 : DFQD1BWP7T port map(CP => clk, D => n_57, Q => bit_counter(3));
  g90196 : CKND2D0BWP7T port map(A1 => n_158, A2 => n_489, ZN => n_405);
  MOSI_shift_reg_14 : DFQD1BWP7T port map(CP => clk, D => n_63, Q => MOSI_shift(14));
  state_reg_1 : DFQD1BWP7T port map(CP => clk, D => n_64, Q => state(1));
  g90180 : INVD1BWP7T port map(I => n_751, ZN => n_749);
  g90205 : NR2D1BWP7T port map(A1 => n_578, A2 => n_105, ZN => n_272);
  g90207 : ND2D1BWP7T port map(A1 => n_158, A2 => MOSI_shift(3), ZN => n_771);
  g90073 : NR2XD0BWP7T port map(A1 => n_135, A2 => n_662, ZN => n_115);
  g90148 : OAI21D0BWP7T port map(A1 => n_171, A2 => n_113, B => full_map_14_1(0), ZN => n_114);
  g90140 : OAI21D0BWP7T port map(A1 => n_171, A2 => n_111, B => full_map_14_3(0), ZN => n_112);
  g90138 : OAI21D0BWP7T port map(A1 => n_1260, A2 => n_219, B => full_map_14_8(0), ZN => n_110);
  g90184 : ND2D1BWP7T port map(A1 => n_451, A2 => full_map_14_9(0), ZN => n_109);
  g90147 : OAI21D0BWP7T port map(A1 => n_202, A2 => n_113, B => full_map_14_13(0), ZN => n_108);
  g90225 : MOAI22D0BWP7T port map(A1 => n_106, A2 => n_105, B1 => n_104, B2 => MOSI_shift(4), ZN => n_107);
  g90136 : OAI21D0BWP7T port map(A1 => n_1260, A2 => n_113, B => full_map_14_9(0), ZN => n_103);
  g90267 : INR3D0BWP7T port map(A1 => n_70, B1 => bit_counter(2), B2 => n_106, ZN => n_102);
  g90183 : CKND2D0BWP7T port map(A1 => n_451, A2 => full_map_7_10(0), ZN => n_101);
  g90182 : OAI31D0BWP7T port map(A1 => n_9, A2 => n_99, A3 => n_104, B => bit_counter(1), ZN => n_100);
  g89988 : OAI31D0BWP7T port map(A1 => n_844, A2 => n_386, A3 => n_169, B => full_map_5_6(0), ZN => n_98);
  g90028 : OAI31D0BWP7T port map(A1 => n_1010, A2 => n_567, A3 => n_171, B => full_map_2_1(2), ZN => n_97);
  g90187 : INR2D1BWP7T port map(A1 => n_285, B1 => n_202, ZN => n_96);
  g90075 : NR2XD0BWP7T port map(A1 => n_135, A2 => n_446, ZN => n_95);
  g90076 : NR2XD0BWP7T port map(A1 => n_116, A2 => n_446, ZN => n_94);
  g90227 : MOAI22D0BWP7T port map(A1 => n_78, A2 => n_637, B1 => n_1150, B2 => MOSI_shift(4), ZN => n_93);
  g90132 : OAI21D0BWP7T port map(A1 => n_1260, A2 => n_111, B => full_map_14_11(0), ZN => n_92);
  g90077 : NR2XD0BWP7T port map(A1 => n_135, A2 => n_485, ZN => n_91);
  g90130 : OAI21D0BWP7T port map(A1 => n_1260, A2 => n_89, B => full_map_14_10(0), ZN => n_90);
  g90219 : OA22D0BWP7T port map(A1 => n_464, A2 => n_252, B1 => n_0, B2 => n_439, Z => n_88);
  g90135 : OAI21D0BWP7T port map(A1 => n_1260, A2 => n_86, B => full_map_10_8(0), ZN => n_87);
  g90195 : CKND2D1BWP7T port map(A1 => n_354, A2 => n_85, ZN => n_632);
  g90197 : NR2D1BWP7T port map(A1 => n_343, A2 => n_628, ZN => n_640);
  g90200 : IND2D1BWP7T port map(A1 => n_84, B1 => MOSI_shift(6), ZN => n_1236);
  g90206 : ND2D1BWP7T port map(A1 => n_354, A2 => n_105, ZN => n_751);
  g90152 : OAI21D0BWP7T port map(A1 => n_169, A2 => n_219, B => full_map_14_4(0), ZN => n_83);
  g90154 : OAI21D0BWP7T port map(A1 => n_169, A2 => n_111, B => full_map_14_7(0), ZN => n_82);
  g90155 : OAI21D0BWP7T port map(A1 => n_169, A2 => n_89, B => full_map_14_6(0), ZN => n_81);
  g90156 : OAI21D0BWP7T port map(A1 => n_169, A2 => n_113, B => full_map_14_5(0), ZN => n_80);
  g90209 : OAI22D0BWP7T port map(A1 => n_78, A2 => n_367, B1 => n_106, B2 => n_909, ZN => n_79);
  g90212 : OAI22D0BWP7T port map(A1 => n_78, A2 => n_76, B1 => n_106, B2 => n_596, ZN => n_77);
  g90186 : INR2D1BWP7T port map(A1 => n_285, B1 => n_171, ZN => n_75);
  g90213 : OAI22D0BWP7T port map(A1 => n_78, A2 => n_105, B1 => n_106, B2 => n_367, ZN => n_74);
  g90228 : MOAI22D0BWP7T port map(A1 => n_78, A2 => n_909, B1 => n_1150, B2 => MOSI_shift(0), ZN => n_73);
  g90226 : MOAI22D0BWP7T port map(A1 => n_106, A2 => n_76, B1 => n_104, B2 => MOSI_shift(9), ZN => n_72);
  g90220 : MOAI22D0BWP7T port map(A1 => n_106, A2 => bit_counter(0), B1 => n_99, B2 => n_70, ZN => n_71);
  g90216 : MOAI22D0BWP7T port map(A1 => n_106, A2 => n_637, B1 => n_104, B2 => MOSI_shift(6), ZN => n_69);
  g90214 : OAI22D0BWP7T port map(A1 => n_78, A2 => n_596, B1 => n_106, B2 => n_16, ZN => n_68);
  g90168 : MOAI22D0BWP7T port map(A1 => n_391, A2 => n_10, B1 => n_118, B2 => n_519, ZN => n_159);
  g90169 : MAOI22D0BWP7T port map(A1 => n_118, A2 => n_1080, B1 => n_634, B2 => n_844, ZN => n_826);
  g90229 : AOI21D0BWP7T port map(A1 => n_30, A2 => full_map_2_0(0), B => n_512, ZN => n_294);
  g90167 : MOAI22D0BWP7T port map(A1 => n_391, A2 => n_366, B1 => n_118, B2 => n_67, ZN => n_160);
  g90264 : INVD0BWP7T port map(I => n_589, ZN => n_225);
  g90191 : NR2D1BWP7T port map(A1 => n_343, A2 => n_662, ZN => n_478);
  g90193 : ND2D1BWP7T port map(A1 => n_354, A2 => full_map_1_2(0), ZN => n_793);
  g90238 : CKND1BWP7T port map(I => n_896, ZN => n_601);
  g90198 : NR2D1BWP7T port map(A1 => n_343, A2 => n_367, ZN => n_240);
  g90242 : CKND1BWP7T port map(I => n_827, ZN => n_804);
  g90203 : IND2D1BWP7T port map(A1 => n_84, B1 => n_519, ZN => n_1232);
  g90202 : OR2D1BWP7T port map(A1 => n_1203, A2 => MOSI_shift(5), Z => n_1242);
  g90204 : NR2D1BWP7T port map(A1 => n_343, A2 => MOSI_shift(3), ZN => n_271);
  g90233 : OR2D1BWP7T port map(A1 => n_48, A2 => n_66, Z => n_1022);
  g90222 : AO22D0BWP7T port map(A1 => n_104, A2 => MOSI_shift(11), B1 => MOSI_shift(10), B2 => n_1150, Z => n_65);
  g90033 : AO22D0BWP7T port map(A1 => n_26, A2 => n_66, B1 => n_12, B2 => n_21, Z => n_64);
  g90224 : AO22D0BWP7T port map(A1 => n_104, A2 => MOSI_shift(14), B1 => MOSI_shift(13), B2 => n_1150, Z => n_63);
  g90159 : NR3D0BWP7T port map(A1 => n_171, A2 => n_781, A3 => n_416, ZN => n_62);
  g90218 : AO22D0BWP7T port map(A1 => n_104, A2 => MOSI_shift(13), B1 => MOSI_shift(12), B2 => n_1150, Z => n_61);
  g90164 : OAI22D0BWP7T port map(A1 => n_391, A2 => n_711, B1 => n_419, B2 => n_366, ZN => n_454);
  g90272 : AOI21D0BWP7T port map(A1 => n_1015, A2 => full_map_2_1(2), B => n_60, ZN => n_851);
  g90232 : ND2D1BWP7T port map(A1 => n_55, A2 => n_1146, ZN => n_208);
  g90239 : INVD1BWP7T port map(I => n_343, ZN => n_158);
  g90257 : ND2D1BWP7T port map(A1 => n_523, A2 => n_967, ZN => n_896);
  g90261 : ND2D1BWP7T port map(A1 => n_523, A2 => n_1087, ZN => n_827);
  g90223 : AO22D0BWP7T port map(A1 => n_104, A2 => MOSI_shift(10), B1 => MOSI_shift(9), B2 => n_1150, Z => n_59);
  g90271 : OAI21D0BWP7T port map(A1 => n_70, A2 => n_17, B => n_78, ZN => n_58);
  g90217 : AO32D1BWP7T port map(A1 => n_1150, A2 => n_70, A3 => bit_counter(2), B1 => n_324, B2 => bit_counter(3), Z => n_57);
  g90208 : AO22D0BWP7T port map(A1 => n_104, A2 => MOSI_shift(12), B1 => MOSI_shift(11), B2 => n_1150, Z => n_56);
  g90235 : INVD0BWP7T port map(I => n_512, ZN => n_388);
  g90240 : CKND1BWP7T port map(I => n_354, ZN => n_578);
  g90247 : ND2D1BWP7T port map(A1 => n_523, A2 => n_992, ZN => n_373);
  g90230 : ND2D1BWP7T port map(A1 => n_55, A2 => n_1015, ZN => n_213);
  g90231 : ND2D1BWP7T port map(A1 => n_55, A2 => n_941, ZN => n_197);
  g90234 : CKND1BWP7T port map(I => n_239, ZN => n_348);
  g90282 : ND2D1BWP7T port map(A1 => n_523, A2 => n_1017, ZN => n_589);
  g90178 : INVD1BWP7T port map(I => n_54, ZN => n_182);
  g90248 : ND2D1BWP7T port map(A1 => n_462, A2 => n_1087, ZN => n_279);
  g90307 : INVD0BWP7T port map(I => n_52, ZN => n_53);
  g90145 : OAI21D0BWP7T port map(A1 => n_50, A2 => n_46, B => n_28, ZN => n_51);
  g89917 : NR2D0BWP7T port map(A1 => n_29, A2 => n_47, ZN => n_49);
  g90269 : OAI22D0BWP7T port map(A1 => n_20, A2 => n_47, B1 => n_46, B2 => MOSI_shift(14), ZN => n_48);
  g90268 : AOI22D0BWP7T port map(A1 => n_1086, A2 => full_map_1_1(2), B1 => n_820, B2 => full_map_2_1(2), ZN => n_45);
  g90201 : NR2XD0BWP7T port map(A1 => n_171, A2 => n_1013, ZN => n_54);
  g90262 : INVD0BWP7T port map(I => n_44, ZN => n_618);
  g90192 : ND2D1BWP7T port map(A1 => n_43, A2 => n_1146, ZN => n_116);
  g90274 : AOI221D0BWP7T port map(A1 => n_596, A2 => full_map_8_0(0), B1 => n_76, B2 => full_map_4_0(0), C => n_39, ZN => n_604);
  g90246 : NR2D0BWP7T port map(A1 => n_628, A2 => n_965, ZN => n_285);
  g90266 : INVD1BWP7T port map(I => n_427, ZN => n_916);
  g90199 : ND2D1BWP7T port map(A1 => n_43, A2 => n_1080, ZN => n_135);
  g90258 : IND2D1BWP7T port map(A1 => n_42, B1 => MOSI_shift(4), ZN => n_343);
  g90270 : AOI22D0BWP7T port map(A1 => n_1086, A2 => full_map_8_4(0), B1 => n_1090, B2 => full_map_11_4(0), ZN => n_41);
  g90318 : CKND2D1BWP7T port map(A1 => n_85, A2 => n_1090, ZN => n_129);
  g90250 : NR2D1BWP7T port map(A1 => n_628, A2 => n_901, ZN => n_239);
  g90265 : INVD0BWP7T port map(I => n_500, ZN => n_437);
  g90190 : ND2D1BWP7T port map(A1 => n_43, A2 => n_941, ZN => n_142);
  g90245 : OR2D1BWP7T port map(A1 => n_42, A2 => n_365, Z => n_84);
  g90194 : ND2D1BWP7T port map(A1 => n_43, A2 => n_1015, ZN => n_148);
  g90288 : INVD1BWP7T port map(I => n_523, ZN => n_774);
  g90281 : AOI221D0BWP7T port map(A1 => n_268, A2 => full_map_4_0(0), B1 => n_40, B2 => full_map_8_0(0), C => n_39, ZN => n_548);
  g90249 : IND2D1BWP7T port map(A1 => n_42, B1 => n_38, ZN => n_1203);
  g90252 : NR2D1BWP7T port map(A1 => n_42, A2 => n_105, ZN => n_451);
  g90251 : NR2D1BWP7T port map(A1 => n_42, A2 => MOSI_shift(3), ZN => n_353);
  g90253 : ND2D1BWP7T port map(A1 => n_634, A2 => n_37, ZN => n_512);
  g90259 : NR2D1BWP7T port map(A1 => n_42, A2 => MOSI_shift(4), ZN => n_354);
  g90243 : IND2D1BWP7T port map(A1 => n_464, B1 => full_map_14_2(0), ZN => n_36);
  g90276 : OAI21D0BWP7T port map(A1 => n_965, A2 => n_222, B => n_390, ZN => n_44);
  g90275 : OAI21D0BWP7T port map(A1 => MOSI_shift(7), A2 => full_map_6_0(0), B => n_15, ZN => n_514);
  g90289 : INVD1BWP7T port map(I => n_628, ZN => n_462);
  g90273 : OAI21D0BWP7T port map(A1 => n_965, A2 => n_679, B => n_390, ZN => n_675);
  g90297 : ND2D1BWP7T port map(A1 => n_1090, A2 => MOSI_shift(8), ZN => n_439);
  g90308 : INVD1BWP7T port map(I => n_337, ZN => n_111);
  g90285 : AOI21D0BWP7T port map(A1 => n_458, A2 => full_map_12_14(0), B => n_35, ZN => n_427);
  g90283 : IOA21D1BWP7T port map(A1 => n_458, A2 => full_map_13_14(0), B => n_34, ZN => n_500);
  g90290 : CKND1BWP7T port map(I => n_104, ZN => n_78);
  g90291 : INVD1BWP7T port map(I => n_1150, ZN => n_106);
  g90293 : NR2XD0BWP7T port map(A1 => n_1013, A2 => n_496, ZN => n_60);
  g90263 : INVD0BWP7T port map(I => n_831, ZN => n_452);
  g90319 : ND2D1BWP7T port map(A1 => n_385, A2 => n_1080, ZN => n_86);
  g90314 : OAI21D0BWP7T port map(A1 => n_901, A2 => n_309, B => n_32, ZN => n_52);
  g90296 : ND2D1BWP7T port map(A1 => n_1080, A2 => n_31, ZN => n_89);
  g90241 : CKND1BWP7T port map(I => n_171, ZN => n_55);
  g90298 : ND2D1BWP7T port map(A1 => n_1080, A2 => n_629, ZN => n_219);
  g90299 : ND2D1BWP7T port map(A1 => n_385, A2 => full_map_10_11(0), ZN => n_468);
  g90279 : IOA21D1BWP7T port map(A1 => n_30, A2 => full_map_3_0(0), B => n_801, ZN => n_118);
  g90301 : ND2D1BWP7T port map(A1 => n_1092, A2 => n_629, ZN => n_113);
  g90236 : INVD1BWP7T port map(I => n_43, ZN => n_202);
  g90303 : NR2XD0BWP7T port map(A1 => n_333, A2 => MOSI_shift(2), ZN => n_523);
  g90141 : AOI211XD0BWP7T port map(A1 => n_25, A2 => state(0), B => state(1), C => SS, ZN => n_29);
  g90360 : INVD1BWP7T port map(I => n_567, ZN => n_85);
  g90324 : NR2XD0BWP7T port map(A1 => n_1010, A2 => n_662, ZN => n_337);
  g90359 : INVD0BWP7T port map(I => n_446, ZN => n_489);
  g90277 : AOI222D0BWP7T port map(A1 => n_458, A2 => full_map_10_14(0), B1 => n_596, B2 => full_map_6_14(0), C1 => n_76, C2 => full_map_2_14(0), ZN => n_603);
  g90278 : AOI222D0BWP7T port map(A1 => n_458, A2 => full_map_11_0(0), B1 => n_596, B2 => full_map_7_0(0), C1 => n_76, C2 => full_map_3_0(0), ZN => n_419);
  g90254 : NR2XD0BWP7T port map(A1 => n_18, A2 => n_105, ZN => n_43);
  g90280 : AOI222D0BWP7T port map(A1 => n_458, A2 => full_map_11_14(0), B1 => n_596, B2 => full_map_7_14(0), C1 => n_76, C2 => full_map_3_14(0), ZN => n_831);
  g90284 : AOI222D0BWP7T port map(A1 => n_458, A2 => full_map_13_0(0), B1 => n_40, B2 => full_map_9_0(0), C1 => n_268, C2 => full_map_5_0(0), ZN => n_391);
  g90304 : ND2D1BWP7T port map(A1 => n_38, A2 => MOSI_shift(2), ZN => n_628);
  g90305 : ND2D1BWP7T port map(A1 => n_28, A2 => n_46, ZN => n_104);
  g90256 : ND2D1BWP7T port map(A1 => n_22, A2 => MOSI_shift(3), ZN => n_169);
  g90332 : INVD1BWP7T port map(I => n_833, ZN => n_1015);
  g90287 : INVD0BWP7T port map(I => n_401, ZN => n_27);
  g90215 : OAI21D0BWP7T port map(A1 => n_25, A2 => SS, B => n_4, ZN => n_26);
  g90317 : AOI22D0BWP7T port map(A1 => n_1087, A2 => full_map_0_0(0), B1 => n_1017, B2 => full_map_1_0(0), ZN => n_557);
  g90315 : OAI21D0BWP7T port map(A1 => n_893, A2 => n_222, B => n_710, ZN => n_755);
  g90311 : INVD0BWP7T port map(I => n_708, ZN => n_555);
  g90309 : INVD0BWP7T port map(I => n_801, ZN => n_460);
  g90310 : INVD1BWP7T port map(I => n_598, ZN => n_551);
  g90323 : MAOI22D0BWP7T port map(A1 => n_40, A2 => full_map_10_0(0), B1 => n_24, B2 => full_map_6_0(0), ZN => n_634);
  g90302 : IND2D1BWP7T port map(A1 => n_23, B1 => MOSI_shift(14), ZN => n_42);
  g90362 : INVD1BWP7T port map(I => n_385, ZN => n_487);
  g90331 : INVD1BWP7T port map(I => n_1086, ZN => n_781);
  g90363 : CKND1BWP7T port map(I => n_629, ZN => n_485);
  g90260 : ND2D1BWP7T port map(A1 => n_22, A2 => n_105, ZN => n_171);
  g90306 : AN2D1BWP7T port map(A1 => n_21, A2 => n_47, Z => n_1150);
  g90329 : CKND1BWP7T port map(I => n_21, ZN => n_20);
  g90364 : INVD0BWP7T port map(I => n_662, ZN => n_31);
  g90316 : AO22D0BWP7T port map(A1 => n_268, A2 => full_map_4_14(0), B1 => full_map_8_14(0), B2 => n_40, Z => n_35);
  g90338 : ND2D0BWP7T port map(A1 => n_1087, A2 => full_map_1_14(0), ZN => n_32);
  g90313 : AOI22D0BWP7T port map(A1 => n_268, A2 => full_map_5_14(0), B1 => n_40, B2 => full_map_9_14(0), ZN => n_34);
  g90378 : INR3D0BWP7T port map(A1 => bit_counter(3), B1 => n_6, B2 => n_17, ZN => n_99);
  g90321 : AOI22D0BWP7T port map(A1 => n_268, A2 => full_map_8_0(0), B1 => n_40, B2 => full_map_12_0(0), ZN => n_558);
  g90330 : INVD1BWP7T port map(I => n_38, ZN => n_333);
  g90350 : ND2D1BWP7T port map(A1 => n_1087, A2 => full_map_1_0(0), ZN => n_664);
  g90361 : INVD1BWP7T port map(I => n_416, ZN => n_422);
  g90325 : AOI22D0BWP7T port map(A1 => n_268, A2 => full_map_7_0(0), B1 => n_40, B2 => full_map_11_0(0), ZN => n_801);
  g90384 : NR2D1BWP7T port map(A1 => n_417, A2 => MOSI_shift(2), ZN => n_385);
  g90366 : INVD1BWP7T port map(I => n_941, ZN => n_844);
  g90354 : ND2D1BWP7T port map(A1 => n_1087, A2 => n_16, ZN => n_833);
  g90353 : NR2XD0BWP7T port map(A1 => n_901, A2 => MOSI_shift(6), ZN => n_1086);
  g90367 : INVD1BWP7T port map(I => n_1117, ZN => n_1090);
  g90312 : AOI22D0BWP7T port map(A1 => n_458, A2 => full_map_10_0(0), B1 => n_76, B2 => full_map_2_0(0), ZN => n_15);
  g90328 : INVD0BWP7T port map(I => n_651, ZN => n_14);
  g90358 : INVD0BWP7T port map(I => n_412, ZN => n_13);
  g90339 : INR2D0BWP7T port map(A1 => full_map_12_0(0), B1 => n_365, ZN => n_39);
  g90244 : AN2D0BWP7T port map(A1 => n_25, A2 => n_12, Z => n_50);
  g90295 : ND2D1BWP7T port map(A1 => n_1146, A2 => MOSI_shift(7), ZN => n_401);
  g90349 : NR2D1BWP7T port map(A1 => n_985, A2 => n_538, ZN => n_526);
  g90322 : AOI22D0BWP7T port map(A1 => n_967, A2 => full_map_0_14(0), B1 => n_992, B2 => full_map_1_14(0), ZN => n_390);
  g90326 : AOI22D0BWP7T port map(A1 => n_268, A2 => full_map_7_14(0), B1 => n_40, B2 => full_map_11_14(0), ZN => n_598);
  g90348 : ND2D1BWP7T port map(A1 => n_1087, A2 => full_map_1_2(0), ZN => n_704);
  g90300 : ND2D1BWP7T port map(A1 => n_1146, A2 => MOSI_shift(8), ZN => n_464);
  g90385 : NR2D1BWP7T port map(A1 => n_365, A2 => MOSI_shift(2), ZN => n_629);
  g90327 : AOI22D0BWP7T port map(A1 => n_268, A2 => full_map_6_14(0), B1 => n_40, B2 => full_map_10_14(0), ZN => n_708);
  g90365 : INVD1BWP7T port map(I => n_820, ZN => n_1009);
  g90381 : ND2D1BWP7T port map(A1 => n_30, A2 => MOSI_shift(2), ZN => n_446);
  g90382 : ND2D1BWP7T port map(A1 => n_30, A2 => n_367, ZN => n_567);
  g90333 : INVD1BWP7T port map(I => n_1010, ZN => n_1092);
  g90334 : INVD1BWP7T port map(I => n_1080, ZN => n_1013);
  g90337 : CKND2D0BWP7T port map(A1 => n_40, A2 => full_map_10_12(0), ZN => n_11);
  g90294 : IND2D1BWP7T port map(A1 => n_8, B1 => MOSI_shift(4), ZN => n_18);
  g90341 : ND2D1BWP7T port map(A1 => n_458, A2 => full_map_14_0(0), ZN => n_37);
  g90345 : NR2D1BWP7T port map(A1 => n_17, A2 => state(0), ZN => n_21);
  g90352 : NR2D1BWP7T port map(A1 => n_455, A2 => MOSI_shift(6), ZN => n_38);
  g90351 : ND2D1BWP7T port map(A1 => n_967, A2 => full_map_1_14(0), ZN => n_710);
  g90383 : ND2D1BWP7T port map(A1 => n_268, A2 => n_367, ZN => n_416);
  g90379 : ND2D1BWP7T port map(A1 => n_40, A2 => MOSI_shift(2), ZN => n_412);
  g90386 : ND2D1BWP7T port map(A1 => n_458, A2 => MOSI_shift(2), ZN => n_662);
  g90388 : NR2D1BWP7T port map(A1 => n_10, A2 => MOSI_shift(1), ZN => n_941);
  g90356 : NR2D1BWP7T port map(A1 => n_893, A2 => n_16, ZN => n_1080);
  g90355 : ND2D1BWP7T port map(A1 => n_967, A2 => MOSI_shift(6), ZN => n_1010);
  g90336 : NR2D0BWP7T port map(A1 => n_17, A2 => bit_counter(0), ZN => n_9);
  g90342 : IND2D1BWP7T port map(A1 => n_17, B1 => state(0), ZN => n_23);
  g90292 : NR2XD0BWP7T port map(A1 => n_8, A2 => MOSI_shift(4), ZN => n_22);
  g90340 : OR2D1BWP7T port map(A1 => n_17, A2 => n_47, Z => n_28);
  g90377 : AOI21D0BWP7T port map(A1 => MOSI_shift(5), A2 => full_map_2_0(0), B => n_670, ZN => n_672);
  g90343 : ND2D1BWP7T port map(A1 => n_967, A2 => full_map_1_2(0), ZN => n_651);
  g90347 : ND2D1BWP7T port map(A1 => n_40, A2 => full_map_8_12(0), ZN => n_616);
  g90346 : NR2D1BWP7T port map(A1 => n_46, A2 => state(1), ZN => n_66);
  g90344 : ND2D1BWP7T port map(A1 => n_967, A2 => full_map_1_13(1), ZN => n_621);
  g90380 : ND2D1BWP7T port map(A1 => n_268, A2 => MOSI_shift(2), ZN => n_386);
  g90387 : NR2D1BWP7T port map(A1 => n_10, A2 => n_909, ZN => n_820);
  g90335 : INVD1BWP7T port map(I => n_1146, ZN => n_1052);
  g90389 : ND2D1BWP7T port map(A1 => n_519, A2 => MOSI_shift(1), ZN => n_1117);
  g90369 : AOI22D0BWP7T port map(A1 => n_76, A2 => full_map_2_2(0), B1 => n_596, B2 => full_map_6_2(0), ZN => n_382);
  g90408 : INVD0BWP7T port map(I => n_268, ZN => n_24);
  g90405 : INVD0BWP7T port map(I => n_10, ZN => n_269);
  g90320 : IND4D0BWP7T port map(A1 => bit_counter(1), B1 => bit_counter(3), B2 => n_7, B3 => n_6, ZN => n_25);
  g90406 : CKND1BWP7T port map(I => n_67, ZN => n_711);
  g90412 : INVD1BWP7T port map(I => n_965, ZN => n_1017);
  g90411 : CKND1BWP7T port map(I => n_992, ZN => n_985);
  g90414 : INVD1BWP7T port map(I => n_893, ZN => n_1087);
  g90368 : INVD0BWP7T port map(I => n_324, ZN => n_5);
  g90393 : INVD0BWP7T port map(I => n_366, ZN => n_513);
  g90373 : AOI22D0BWP7T port map(A1 => n_637, A2 => full_map_0_0(0), B1 => MOSI_shift(5), B2 => full_map_1_0(0), ZN => n_666);
  g90392 : INVD0BWP7T port map(I => n_336, ZN => n_345);
  g90407 : INVD1BWP7T port map(I => n_455, ZN => n_30);
  g90409 : INVD1BWP7T port map(I => n_40, ZN => n_417);
  g90410 : CKND1BWP7T port map(I => n_458, ZN => n_365);
  g90413 : INVD1BWP7T port map(I => n_967, ZN => n_901);
  g90357 : NR2XD0BWP7T port map(A1 => n_798, A2 => MOSI_shift(1), ZN => n_1146);
  g90372 : IND3D1BWP7T port map(A1 => MOSI_shift(14), B1 => state(1), B2 => state(0), ZN => n_8);
  g90376 : AOI22D0BWP7T port map(A1 => MOSI_shift(8), A2 => full_map_12_14(0), B1 => MOSI_shift(7), B2 => full_map_8_14(0), ZN => n_550);
  g90417 : NR2D1BWP7T port map(A1 => n_16, A2 => MOSI_shift(5), ZN => n_67);
  g90397 : NR2D1BWP7T port map(A1 => MOSI_shift(5), A2 => n_287, ZN => n_670);
  g90401 : ND2D1BWP7T port map(A1 => n_76, A2 => full_map_3_2(1), ZN => n_336);
  g90374 : AOI22D0BWP7T port map(A1 => MOSI_shift(8), A2 => full_map_13_0(0), B1 => MOSI_shift(7), B2 => full_map_9_0(0), ZN => n_492);
  g90416 : CKND2D1BWP7T port map(A1 => MOSI_shift(5), A2 => n_16, ZN => n_10);
  g90399 : INR2D1BWP7T port map(A1 => bit_counter(1), B1 => n_7, ZN => n_70);
  g90403 : ND2D1BWP7T port map(A1 => n_637, A2 => n_16, ZN => n_366);
  g90422 : NR2D1BWP7T port map(A1 => n_637, A2 => n_909, ZN => n_992);
  g90421 : NR2D1BWP7T port map(A1 => n_76, A2 => n_596, ZN => n_458);
  g90420 : NR2D1BWP7T port map(A1 => n_76, A2 => MOSI_shift(7), ZN => n_40);
  g90424 : NR2XD0BWP7T port map(A1 => n_909, A2 => MOSI_shift(5), ZN => n_967);
  g90391 : INVD0BWP7T port map(I => n_12, ZN => n_4);
  g90370 : AOI22D0BWP7T port map(A1 => MOSI_shift(8), A2 => full_map_13_14(0), B1 => MOSI_shift(7), B2 => full_map_9_14(0), ZN => n_554);
  g90371 : AOI22D0BWP7T port map(A1 => MOSI_shift(8), A2 => full_map_14_0(0), B1 => MOSI_shift(7), B2 => full_map_10_0(0), ZN => n_466);
  g90415 : ND2D1BWP7T port map(A1 => n_367, A2 => n_76, ZN => n_334);
  g90375 : AOI22D0BWP7T port map(A1 => MOSI_shift(8), A2 => full_map_12_0(0), B1 => MOSI_shift(7), B2 => full_map_8_0(0), ZN => n_418);
  g90400 : ND2D1BWP7T port map(A1 => state(0), A2 => n_3, ZN => n_46);
  g90394 : INVD1BWP7T port map(I => n_798, ZN => n_519);
  g90402 : ND2D1BWP7T port map(A1 => state(1), A2 => n_3, ZN => n_17);
  g90418 : CKND2D1BWP7T port map(A1 => n_596, A2 => n_76, ZN => n_455);
  g90419 : NR2D1BWP7T port map(A1 => n_596, A2 => MOSI_shift(8), ZN => n_268);
  g90423 : ND2D1BWP7T port map(A1 => n_909, A2 => MOSI_shift(5), ZN => n_965);
  g90425 : ND2D1BWP7T port map(A1 => n_637, A2 => n_909, ZN => n_893);
  g90390 : OA21D1BWP7T port map(A1 => state(0), A2 => state(1), B => n_3, Z => n_324);
  g90396 : INR2D1BWP7T port map(A1 => full_map_0_0(0), B1 => MOSI_shift(1), ZN => n_493);
  g90404 : ND2D1BWP7T port map(A1 => MOSI_shift(5), A2 => MOSI_shift(6), ZN => n_798);
  g90395 : INR2XD0BWP7T port map(A1 => SCLK, B1 => SS, ZN => n_12);
  g90398 : NR2XD0BWP7T port map(A1 => SS, A2 => SCLK, ZN => n_47);
  g90426 : INVD1BWP7T port map(I => reset, ZN => n_3);
  drc_bufs90628 : INVD4BWP7T port map(I => n_1252, ZN => MISO);
  full_map_reg_14_1_0 : DFD1BWP7T port map(CP => clk, D => n_194, Q => full_map_14_1(0), QN => n_2);
  full_map_reg_5_2_0 : DFD1BWP7T port map(CP => clk, D => n_317, Q => full_map_5_2(0), QN => n_316);
  full_map_reg_3_14_0 : DFD1BWP7T port map(CP => clk, D => n_264, Q => full_map_3_14(0), QN => n_263);
  full_map_reg_1_14_0 : DFD1BWP7T port map(CP => clk, D => n_245, Q => full_map_1_14(0), QN => n_244);
  full_map_reg_11_4_0 : DFD1BWP7T port map(CP => clk, D => n_302, Q => full_map_11_4(0), QN => n_301);
  full_map_reg_2_14_0 : DFD1BWP7T port map(CP => clk, D => n_261, Q => full_map_2_14(0), QN => n_432);
  full_map_reg_6_2_0 : DFD1BWP7T port map(CP => clk, D => n_318, Q => full_map_6_2(0), QN => n_411);
  full_map_reg_1_13_1 : DFD1BWP7T port map(CP => clk, D => n_278, Q => full_map_1_13(1), QN => n_222);
  full_map_reg_14_14_0 : DFD1BWP7T port map(CP => clk, D => n_251, Q => full_map_14_14(0), QN => n_465);
  full_map_reg_1_1_2 : DFD1BWP7T port map(CP => clk, D => n_312, Q => full_map_1_1(2), QN => n_570);
  full_map_reg_1_2_0 : DFD1BWP7T port map(CP => clk, D => n_246, Q => full_map_1_2(0), QN => n_538);
  MOSI_shift_reg_6 : DFD1BWP7T port map(CP => clk, D => n_69, Q => MOSI_shift(6), QN => n_16);
  full_map_reg_4_2_0 : DFD1BWP7T port map(CP => clk, D => n_314, Q => full_map_4_2(0), QN => n_546);
  MOSI_shift_reg_5 : DFD1BWP7T port map(CP => clk, D => n_93, Q => MOSI_shift(5), QN => n_637);
  MOSI_shift_reg_7 : DFD1BWP7T port map(CP => clk, D => n_68, Q => MOSI_shift(7), QN => n_596);
  full_map_reg_8_12_0 : DFD1BWP7T port map(CP => clk, D => n_250, Q => full_map_8_12(0), QN => n_1);
  full_map_reg_14_13_0 : DFD1BWP7T port map(CP => clk, D => n_188, Q => full_map_14_13(0), QN => n_0);
  full_map_reg_0_14_0 : DFD1BWP7T port map(CP => clk, D => n_305, Q => full_map_0_14(0), QN => n_304);
  bit_counter_reg_2 : DFD1BWP7T port map(CP => clk, D => n_242, Q => bit_counter(2), QN => n_6);
  full_map_reg_1_0_0 : DFD1BWP7T port map(CP => clk, D => n_288, Q => full_map_1_0(0), QN => n_287);
  bit_counter_reg_0 : DFD1BWP7T port map(CP => clk, D => n_178, Q => bit_counter(0), QN => n_7);
  full_map_reg_2_2_0 : DFD1BWP7T port map(CP => clk, D => n_315, Q => full_map_2_2(0), QN => n_579);
  full_map_reg_2_0_0 : DFD1BWP7T port map(CP => clk, D => n_310, Q => full_map_2_0(0), QN => n_309);
  full_map_reg_14_12_0 : DFD1BWP7T port map(CP => clk, D => n_253, Q => full_map_14_12(0), QN => n_252);
  full_map_reg_0_1_0 : DFD1BWP7T port map(CP => clk, D => n_284, Q => full_map_0_1(0), QN => n_566);
  full_map_reg_2_1_2 : DFD1BWP7T port map(CP => clk, D => n_206, Q => full_map_2_1(2), QN => n_488);
  full_map_reg_4_1_2 : DFD1BWP7T port map(CP => clk, D => n_199, Q => full_map_4_1(2), QN => n_496);
  full_map_reg_1_13_0 : DFD1BWP7T port map(CP => clk, D => n_381, Q => full_map_1_13(0), QN => n_679);
  MOSI_shift_reg_3 : DFD1BWP7T port map(CP => clk, D => n_74, Q => MOSI_shift(3), QN => n_105);
  MOSI_shift_reg_2 : DFD1BWP7T port map(CP => clk, D => n_79, Q => MOSI_shift(2), QN => n_367);
  MOSI_shift_reg_8 : DFD1BWP7T port map(CP => clk, D => n_77, Q => MOSI_shift(8), QN => n_76);
  MOSI_shift_reg_1 : DFD1BWP7T port map(CP => clk, D => n_73, Q => MOSI_shift(1), QN => n_909);
  MISO_shift_reg_72 : DFD0BWP7T port map(CP => clk, D => n_560, Q => MISO_shift(72), QN => n_1252);
  g2 : IND4D0BWP7T port map(A1 => n_983, B1 => n_1116, B2 => n_1231, B3 => n_1242, ZN => n_1256);
  g90699 : IND4D0BWP7T port map(A1 => n_377, B1 => n_958, B2 => n_1050, B3 => n_846, ZN => n_1257);
  g90700 : IND2D1BWP7T port map(A1 => n_369, B1 => n_804, ZN => n_1258);
  g90701 : IND2D1BWP7T port map(A1 => n_169, B1 => n_385, ZN => n_1259);
  g90702 : IND2D1BWP7T port map(A1 => n_18, B1 => n_105, ZN => n_1260);

end synthesised;
