configuration color_ctrl_behavioural_cfg of color_ctrl is
   for behavioural
   end for;
end color_ctrl_behavioural_cfg;
