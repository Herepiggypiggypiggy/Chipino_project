configuration display_ctrl_behavioural_cfg of display_ctrl is
   for behavioural
   end for;
end display_ctrl_behavioural_cfg;
