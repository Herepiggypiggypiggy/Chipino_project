configuration player_fsm_behaviour_cfg of player_fsm is
   for behaviour
   end for;
end player_fsm_behaviour_cfg;
