entity display_ctrl_tb2 is
end display_ctrl_tb2;

