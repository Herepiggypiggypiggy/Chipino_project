configuration module_test_synthesised_cfg of module_test is
   for synthesised
   end for;
end module_test_synthesised_cfg;
