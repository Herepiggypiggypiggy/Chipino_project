configuration stable_map_behaviour_cfg of stable_map is
   for behaviour
   end for;
end stable_map_behaviour_cfg;
