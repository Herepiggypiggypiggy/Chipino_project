configuration spi_v3_behaviour_cfg of spi_v3 is
   for behaviour
   end for;
end spi_v3_behaviour_cfg;
