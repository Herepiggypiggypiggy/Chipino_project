entity display_ctrl_tb is
end display_ctrl_tb;

